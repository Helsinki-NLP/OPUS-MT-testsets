Ии.
Гыт микигыт?
Гымнин нынны Том.
