Beskrivning:  
I samband med skrivandet av Byggðasögu Skagafjarðar, Skagafjörðurs bygdehistoria, har en omfattande undersökning genomförts av forntida ödemark i dalarna och på hedarna i Skagafjörður. 
I samarbete med Hjalti Pálsson, historiker och författare av bygdehistoria, och Þór Hjaltalín, naturvårdare för Norðurland vestra, åtog sig den arkeologiska avdelningen vid Byggðasafns Skagfirðinga, Skagafjörðurs bygdemuseum, att ta marksnitt i utvalda lämningar. 
Avsikten var att bestämma ålder av och kanske även vem som byggde dem, och i förekommande fall även om de faktiskt är lämningar.  
Náttúrustofa Norðurlands vestra, Västra nordlandets naturdepartement, deltog också i en del av projektet, där dess medarbetare Helgi Páll Jónsson hjälpte till med pyroklasteranalysen när han arbetade med forskning för sin kandidatavhandling "Gjóskulög í Skagafjörður", Pyroklaster i Skagafjörður. 
Dessutom analyserade Magnús Sigurgeirsson pyroklasterprover som togs vid den gamla gården Tunga i Vesturdalur och hans analysrapport bifogas. 
De utvalda platserna hittades av Hjalti Pálsson under hans forskningsresor, men han har sökt efter gårdar och områden som är kända från källor men vars läge har inte varit kända. 
I Árnis och Pálls Jordabok beskrivs gården Fögruhlíð enligt följande: "Fagrahlijd. 
Ödegård framför Nýjabær har varit öde länge, även om det finns synliga byggnationslämningar, staket runt ängen och ruiner. 
Området runt tunet är helt förfallet och svårt att bygga på, eftersom det inte finns någon slåtteräng så pass nära att odling kan upprättas. 
Annars är betesmarkerna här anmärkningsvärt goda både på sommaren och vintern" (Árni Magnússon och Páll Vídalín, 1930: 65). 
Cirka 8,5 km framför Ábær, 350 m.ö.h. och cirka 250 meter framför Hjálmarsselslækur finns två raviner, den yttre är bevuxen och mycket bredare än den södra, till hälften bevuxna, ravinen. 
Mellan dem finns en smal tunga eller sektor, 25-30 meter bred, täckt med buskar. 
Längst ner i denna sektor nere vid stranden av Jökulsá är det otydligt och i nersjunkna i marken finns lämningar av hus och trädgårdsodling. 
Ruinen är gräsbevuxen och det verkar finnas fyra avdelningar på en yta med yttermått på cirka 10x8 m. 
Cirka 10 m utanför (norr om) ruinen finns ett otydligt trädgårdsområde, täckt av jord, delvis gömt under ljung och pilbuskar. 
Trädgårdsområdet ligger ungefär i öst-västlig riktning och är cirka 15 meter långt. 
Det finns en djup grop strax norr om ruinen. 
Jökulsá har eroderat tiotals, om inte hundratals, meter mark och floden har brutit banken hela vägen upp till ruinerna och där är den ungefär 10 meter hög (Hjalti Pálsson, 2007). 
Ruinområdet verkar delvis ha försvunnit framför den eroderade flodbanken.  
Hela området är täckt av buskar och det var inte möjligt att säkert identifiera gärdesgården eller ruinerna. 
Ytterligare beskrivning: 
Den forntida gården Fagrahlíð i Austurdalur i Skagafjörður. 
Fotot är taget mot öster i ett marksnitt, för analys, som tagits längs en vägg i ruinen. 
Beskrivning: 
Den så kallade Herpisgerði ligger långt söder om Hofsá, i princip rakt mittöver Hrafnhóll öster om Hjaltadalsá, några hundra meter öster om floden, men från gården är det cirka hundra meter torvmark upp till bruket. 
Det kan ha legat en gammal gård här. 
Det har funnits en rejäl gärdesgård runtom, mestadels cirkulär, som sjunkit ner i den sydvästra delen av myren, men det finns fortfarande en tydlig odling i marken innanför gärdesgården. 
Man kan anta att markytan på gården är minst 1,5 hektar. 
Huvuddelen av ruinen är lång och mycket förstörd och går i höjd med marken där den står, det verkar ha varit en fårfålla eller kanske ett [avskilt beläget] fårhus tillhörande Hólar, även om ingen gård syns till. 
Den ligger i öst-västlig riktning, dörren vetter åt väster direkt mot Hrafnhóll. 
Total längd, ca 21 m på insidan. 
Från ruinen och till båda sidorna är ruinen över 20 meter lång. 
Förmodligen ett äldre hus. 
Ett tydligt fält ligger öster om ruinerna av [det avskilt belägna] fårhuset. 
Österut under gården, strax söder om den östra änden av ovannämnda ruin, finns en annan lång ruin, mycket äldre och som går i nord-sydlig riktning, även den ungefär 22-23 meter lång på utsidan, uppdelad i tre eller fyra avdelningar, 5-6 meter bred på utsidan. 
Ruinerna är ganska otydliga och det är svårt att avgöra vilken typ av hus dessa har varit. 
Några meter öster om huvudruinen och vallen finns en stor rektangulär ruin, cirka 8x9 m stor, ganska otydlig och det kan inte ha varit ett hus, snarare en fårfålla. 
Det är den överlägset mest otydliga av dessa tre ruiner. 
Alla dessa lämningar är stora, märkliga och svåra att förklara. 
Gårdsbågarna söder om ruinerna är faktiskt tre stycken och i den sydvästra änden av en av dem verkar det finnas små lämningar i marken. 
Ytterligare beskrivning: Herpisgerði - marksnitt 1 i gärdesgården - norra delen Marksnitt 1 - i " gärdesgården " Marksnitt 1 gjordes på östra sidan av gärdesgården. 
Det var 180 cm långt, 60 cm brett och cirka 80 cm djupt. 
Längst ner vid gräsrötterna fanns cirka 0,5 cm tjock svart pyroklaster, H1766. 
Ett orört lager av lössjord [2] ca 10-15 cm tjockt låg omedelbart under gräsrötterna och gick ner till ruinväggen. 
Ruinväggen [4] kan urskiljas längs det längsgående marksnittet, den tjockaste delen i mitten var ca 50 cm hög. 
I marksnitten fanns två detekterbara pyroklasterlager, H1104 och H1300. 
Det fanns mycket lera i ruinen och ovanför väggarna öster om marksnittet fanns ett 10 cm tjockt lager[3] med lera och sand. 
Under ruinväggen fanns ett ungefär lika tjockt rotat grässkikt [5] ungefär 15 cm tjockt. 
Den innehöll rödaktig torvmossa med ett lager av H1104. 
Detta rotade torvlager låg sedan orört direkt ovanpå H1300. 
Under H1300 fanns det ett 10 cm tjockt obearbetat lössjordsskikt ner till H1104 som även det var orört. 
Det fanns inga tecken på en mänsklig boning under H1300.
Tolkning av marksnittet: 
En gärdesgårdsmur har byggts, möjligen på 1300- eller 1400-talet. 
Det var inte möjligt att avgöra om gården hade byggts om och därför kan den ha varit i bruk endast under relativt kort tid. 
Den förföll långt före nedfallet av 1766 års pyroklaster. 
Byggnaden som grävdes ut verkar ha varit ett uthus snarare än en mänsklig boning och verkar ha byggts samtidigt som gärdesgården. 
Byggnaden restes efter år 1300 men förföll och revs långt innan nedfallet av 1766 års pyroklaster.
Beskrivning: 
Nýlendi är en ödegård vars ägor ligger mellan Grindur i Deildardalur i öster och Ennis vid Höfðaströnd i norr. 
Den äldsta noteringen om gården finns i en köpehandling från 1400-talet när marken såldes till biskopssätet i Hólar, då den uppmättes till 25 hundraden (Diplomatarium Islandicum, Íslenskt fornbréfasafn DI IV, s. 553-554). 
I Jordaboken från 1709 är marken för två familjer/gårdar och värderades till 35 hundraden (Árn Magnússons och Pál Vídalíns Jordabok X, s. 244) men 40 hundraden när den såldes av 1802. 
I Johnsens Jordabok från 1847 värderades å andra sidan marken till 36 hundraden (Johnsens Jordabok 1847, s. 270). 
Nu [2013] ägs Nýlendi av Laugabóls ehf (Veðmálabækur Skagafjarðar, Skagafjördurs inteckningsregister, nr. 161/2007). 
Den nuvarande betongbostadsbyggnaden står på Langahóll cirka 60 meter söder om Bæjarhóll, där de övervuxna ruinerna av gården fortfarande är synliga.  
Den gamla gården stod där tills den nuvarande bostadsbyggnaden byggdes 1942. 
Arrende eller avhysning nämns inte i fastighetsregistret från 1709, men två sådana har registrerats i markägarregistret. 
Annars var det lämningar av en namnlös bostadshus, gärdesgård och ruiner som låg i Nýlendishvammur vid Deildardalsá, strax söder om Deildardalsvegur. 
Ingólfur Jónsson, en bonde i Nýlendi, jämnade under sin lantbrukstid både ruinerna och gården med marken med en bulldozer och planerade att odla potatis där, men dessa planer förverkligades aldrig (Svanhildur Guðjónsdóttir, muntlig källa 2013). 
Nýlendiskot heter lämningarna av en gärdesgård med ruinrester cirka 300 m utifrån och upp från gårdshusen i Nýlendi, nära betesmarkerna. 
Det sägs att det varit en bostad där, men inga skriftliga källor stöder dessa berättelser. 
Man tror att det har funnits ett fårhus där, men ortsnamnsregistret innehåller inte tillförlitlig information om stugan. 
Vid Nýlendiskot finns vad som liknar ett övervuxet tun. 
Vid första anblicken finns det en tydlig gärdesgård runt ett igenvuxet tun som mäter 0,7 ha. 
Hö skördades i Nýlendiskot in på 1900-talet, åtminstone fram till 1945 och höet transporterades därifrån på ridhästar sommartid (Svanhildur Guðjónsdóttir, muntlig källa 2013). Vid närmare granskning kan man se att en mycket äldre gärdesgård omger den tidigare nämnda. 
Men den gården har bitvis försvunnit men syns till största delen tydligt, särskilt i norr och öster. 
I söder är den nya gården byggd ovanpå den äldre, som är ganska stor, och det är uppenbart att den inte har byggts runt någon stuga.
En mindre arkeologisk undersökning utfördes av lämningarna vid Nýlendiskot. 
Fyra borrkärneprov togs i den påstådda gårdskullen och dess omgivningar. 
Det visade sig att under ruinerna av fårhusen fanns rester av en gammal bondgård som verkar ha varit i bruk före år 1104. 
Erosionssnittet från den äldre gärdesgården rensades och inspekterades. 
Gärdesgårdsmuren var cirka 60 cm hög och i den fanns torv med mycket H3-pyroklaster men inga bevis för pyroklaster från 1104 eller 1300. 
Ingen pyroklaster kunde detekteras ovanför eller upp längs muren. 
Det var därför inte möjligt att datera den ytterligare, även om det kan anses osannolikt att pyroklastern från 1104 inte skulle finnas i ruinerna om de hade rests efter nedfallet av pyroklastern. 
En mindre erosionsprofil undersöktes även i den yngre trädgården. 
Det var inte möjligt att ytterligare identifiera ruinerna som fanns på gården, men den har byggts ovanpå H1104 pyroklastisk sten. 
Den är dock utan tvekan betydligt yngre med tanke på hur tydlig den är.
Tolkning:
Det har där funnits en gård åtminstone på 1000-talet som förmodligen kom från en bosättning mycket tidigt, ev. redan på 1000-talet. 
Stugan som området är uppkallat efter byggdes efter 1104, troligen mycket senare. 
L-formade ruiner uppe vid den yngre gärdesgården hör antagligen till den. 
Ytterligare beskrivning: 
Stenar på utsidan och väster om en äldre gärdesgård väster om Nýlendiskot. Sett norrut. 
Beskrivning: 
Ödebygd och dalar III. 2008. 
"Gårdshus" i Hólahagi i landet Hólar i Hjaltadalur.
Ett marksnitt togs i en forntida ruin i Hólahagi i trakten av Hólastaður i Hjaltadalur. 
Det finns inga register över gårdar med detta namn (d.v.s. Garðhús) men i närheten av lämningarna finns de så kallade Garðhúsagil och Garðhúsaskriða. 
Det finns tydliga rester av äldre lämningar på platsen, men det finns även rester av någon slags fårfållor, kanske ett senare tiders [avskilt beläget] fårhus. 
Ruinerna ligger längst fram på stranden ovanför och väster om Hjaltadalsá ungefär en kilometer in från Hof och är mycket nedsjunkna i marken. 
Det är en långsträckt ruin som är cirka 20 meter lång och troligen två ruiner eller bihus till väster om den.  
Ovanför dessa ruiner finns två yngre ruiner, möjligen resterna av ett [avskilt beläget] fårhus eller fårfålla. 
Ytterligare beskrivning: 
Utgrävning av ruinerna av en stuga i Hólahagi. 
Sett mot nordväst. 
Marksnitt 1 - taget i den nordvästra kortväggen av en eventuell stugruin Marksnittet togs i den nordvästra kortsidan av den långa ruinen.
En torvvägg hittades, som innehåller fragment av grönaktig pyroklaster, det så kallade bosättningsskiktet, som nedföll 872. 
Det fanns även rikligt med förhistorisk pyroklaster från Hekla i väggen. 
Söder om snittet hade rester av ett svart golvlager förts ner när väggen eller taktorven kollapsat.
Golvskiktet var ett svart fettigt golvskikt, cirka 5-7 cm tjockt med kol, brända ben och gråaktig aska. 
Ovanpå golvskiktet fanns cirka 10 cm orörd tätningsjord och ovanför fanns pyroklasterlager från Hekla från 1104 och 1300. 
Skikten låg upp mot väggen på södersidan och väggen har kollapsat före nedfallet av pyroklastern från 1104. 
Inga pyroklasterskikt hittades längs väggen eller i den kollapsade norra delen av den, annars fanns ett mycket tunt svart pyroklasterskikt strax under gräsrötterna norr om snittet. 
Det kan vara pyroklaster från Hekla som nedföll 1766.
Tolkning av marksnitten:
Detta är ett boningshus, en stuga som troligen har tagits i bruk strax efter det att bosättningsskiktet föll men som revs strax innan pyroklastern från 1104 nedföll. 
Det gick inte att se att det hade funnits en gärdesgård runt byggnaden, men många jordskred har gått i sluttningen runt om och spåren efter gärdesgården och andra byggnationer kan ha försvunnit. 
Beskrivning: 
Bäcken omnämns först i mitten av 1300-talet, men arkeologiska fynd indikerar att området var bebott från de tidigaste bosättningstiderna.
Jordbruket upphörde 1958 och marken är nu en del av Ennis mark och nyttjas därifrån (Byggðasaga Skagafjarðar V, Skagafjörðurs bygdehistoria Volym 5, s. 269-270). 
Inga fler byggnader är uppförda, men gårdskullen är fortfarande tydligt igenkännlig. 
Gärdesgården kan ses delvis till väster och norr om gårdskullen och det finns två ruiner vid dess västra del. 
Cirka 20-50 meter direkt norr om gårdskullen finns otydliga fornlämningar, ruiner av stugor och andra byggnadsrester. 
Borrkärneprov togs i ruiner och gärdesgård, förutom att ett marksnitt togs inne i stugruinerna. 
Ytterligare beskrivning: 
Lækur i Viðvíkursveit. 
Resterna av en fårfålla öster om boningshusruinen. 
Sett söderut.
Beskrivning: 
Den så kallade Herpisgerði ligger långt söder om Hofsá, i princip rakt mittöver Hrafnhóll öster om Hjaltadalsá, några hundra meter öster om floden, men från gården är det cirka hundra meter torvmark upp till bruket. 
Det kan ha legat en gammal gård här. 
Det har funnits en rejäl gärdesgård runtom, mestadels cirkulär, som sjunkit ner i den sydvästra delen av myren, men det finns fortfarande en tydlig odling i marken innanför gärdesgården. 
Man kan anta att markytan på gården är minst 1,5 hektar. 
Huvuddelen av ruinen är lång och mycket förstörd och går i höjd med marken där den står, det verkar ha varit en fårfålla eller kanske ett [avskilt beläget] fårhus tillhörande Hólar, även om ingen gård syns till. 
Den ligger i öst-västlig riktning, dörren vetter åt väster direkt mot Hrafnhóll. 
Total längd, ca 21 m på insidan. 
Från ruinen och till båda sidorna är ruinen över 20 meter lång. 
Förmodligen ett äldre hus. 
Ett tydligt fält ligger öster om ruinerna av [det avskilt belägna] fårhuset. 
Österut under gården, strax söder om den östra änden av ovannämnda ruin, finns en annan lång ruin, mycket äldre och som går i nord-sydlig riktning, även den ungefär 22-23 meter lång på utsidan, uppdelad i tre eller fyra avdelningar, 5-6 meter bred på utsidan. 
Ruinerna är ganska otydliga och det är svårt att avgöra vilken typ av hus dessa har varit. 
Några meter öster om huvudruinen och vallen finns en stor rektangulär ruin, cirka 8x9 m stor, ganska otydlig och det kan inte ha varit ett hus, snarare en fårfålla. 
Det är den överlägset mest otydliga av dessa tre ruiner. 
Alla dessa lämningar är stora, märkliga och svåra att förklara. 
Gårdsbågarna söder om ruinerna är faktiskt tre stycken och i den sydvästra änden av en av dem verkar det finnas små lämningar i marken. 
Ytterligare beskrivning: Herpisgerði - marksnitt 2 i en ruin vid gärdesgård - östra snittet Marksnitt 2 - i en ruin av en stadig gärdesgårdsmur 
Ett annat marksnitt togs sedan i den inre delen av en ruinvägg i en fyrdelad ruin som gränsade till tunet i öster.
Längst ner vid gräsrötterna fanns cirka 0,5 cm tjock svart pyroklaster, H1766. 
Under fanns det cirka 5 cm tjock lössjord [2] ner till ruinväggen. 
Väggen [3] var gjord av torv som innehöll pyroklaster-skiktet Hekla 1300. 
En kollapsad del av torvväggen [4] hittades inne i ruinen men inga tecken på golvskikt hittades.
Tolkning av marksnittet: 
En gärdesgårdsmur har byggts, möjligen på 1300- eller 1400-talet. 
Det var inte möjligt att avgöra om gården hade byggts om och därför kan den ha varit i bruk endast under relativt kort tid. 
Den förföll långt före nedfallet av 1766 års pyroklaster. 
Byggnaden som grävdes ut verkar ha varit ett uthus snarare än en mänsklig boning och verkar ha byggts samtidigt som gärdesgården. 
Byggnaden restes efter år 1300 men förföll och revs långt innan nedfallet av 1766 års pyroklaster.
Beskrivning: 
Marbælisselland ligger precis framför Óslandsselland öster om Seljadalur. 
Den går från Glúmsgil till Strangalæk, och är cirka 2,5 km lång. 
I fastighetsregistret från 1709 står: "Selstaður äger marken i Seljadalur, men har inte användning för avlägsna platser, så andra använder marken i otacksamhet." 
Tyvärr anges inte vem som använder marken i "otacksamhet" eller om andra använder det som fäbodsviste eller endast använder marken för bete. 
Fäbodsruinerna ligger 210 m nedanför Glúmsgil i Seljadalur och där finns tydliga ruiner. 
Huvudruinen är cirka 10x7 m, verkar vara uppdelad i fem bostäder och väggränserna är ganska tydliga. 
Några meter västerut finns fårfållorna, 3x8 m på utsidan, men nära dem verkar det ha funnits ett litet hus, cirka 2x2m. 
Fäboden ligger nära hemmanet vid Glúmsgilslækur och ingår i Óslandsselland och måste ha anlagts där med tillstånd av Óslandsbönderna, såvida inte bäcken har ändrat sitt flöde. 
När Steinar Þórðarson var ung i Háleggstaður fanns det en skyddad del i floden nedanför fäboden som kallades Glúmsgilshylur och det var en av de bästa fiskeplatserna i floden. 
Där finns plana grunder och en vacker fäbod. 
(Byggðasaga Skagafjarðar VII., Skagafjörðurs bygdehistoria volym 7, Hofshreppur, 189) 
Ytterligare beskrivning: 
Marbælissel i Seljadalur. 
Sett österut.
Beskrivning: 
Från början har projektet varit en del av arbetet med att skriva Byggðasagan, Byggdehistoren, nu har fyra framgångsrika volymer publicerats. 
Byggðasagan skiljer sig från andra lokalhistoriska böcker genom att det läggs större vikt vid gårdarnas forntida historia och studiet av alla typer av arkeologiska lämningar som kan läggas till deras historia. 
De två sista volymerna av Byggðasagan innehåller detaljerade kapitel om forntida bosättningar i de inre dalarna i Austurdalur och Vesturdalur, där historien är sammanflätad med resultaten av arkeologiska utgrävningar som har ägt rum på utvalda platser. 
Den forntida gården Risamýr nämns i en forntida källa, men den exakta platsen för gården är okänd. 
I den fjärde volymen av Byggðasögu Skagafjarðar, Skagafjörðurs bygdehistoria, (s. 172-173) finns indikationer på var denna gård sannolikt kan ha legat. 
Området norr om Réttarholt, väster om Héraðsvatn österut under Þormóðsholt, är en enorm sumpmark, våtmark innan gården restes och fram till för en tid sedan, en verklig jättemyr. 
Den forntida brevsamlingen innehåller ett brev om Risamýri från år 1369 då biskop Jón avgör att Hólakirkjas har äganderätt till marken i Risamýr, "i Guds namn, amen." 
Det är oklart om Risamýr var landskapsmark eller ödemark, med det ovan nämnda forntidsbrevet nämner "marken i Risamýr" vilket stöder bilden att Risamýri tidigare var en gård. Vid 1369 var den troligtvis öde för länge sedan och marken låg delvis under Bjarnastaðir och till viss del Flugumýri. 
Ortsnamnet är inte längre känt, men det finns knappast något annat man tänker på än slätmarken nedanför Þormóðsholt och ner till Vötnar. 
Biskopen sa att Risamýri ingick i marken som tillhörde biskopssätet Flugumýr och att den hade nyttjats som sådan i årtionden. 
Får betade där på sommaren och hästar på vintern under mer än 40 år. 
Det verkar som att Risamýri var beläget i Bjarnastaðaland eller att det av vissa ansågs vara en del av den mark som verkar ha ägts av Magnús Grímsson som kanske då bodde i Bjarnastaðir. 
Han fick "ingen invändning i gengäld... till en boning i Bjarnastaðir" och Risamýri tilldömdes sedan till Flugumýri (Fornbréfasafn Íslands III, Islands arkeologiska museum, 252-253). 
Som nämnts i diskussioner runt Bjarnastaðir har det varit en stor mark en gång i tiden, men är det inte längre. 
Det förklaras inte på något annat sätt, så som det verkar, men ursprungligen ingick marken väster om Héraðsvatn. 
Detta har dock inte varit fallet under de senaste århundradena.  
Flugumýri har länge varit känt för att äga marken väster om Þormóðsholt, väster om den nuvarande landsvägen. 
Det bör även noteras att Réttarholts mark ursprungligen var uthyrd under ett arrende från marken i Flugumýr. 
I sin sökning efter "marken Risamýr" har registratorn [Hjalti Pálsson] stannat vid Skiphóll, vilket diskuteras ovan. Den är cirka 60 meter lång, på många ställen ganska stor och bakom den finns gamla ridleder. 
På kullen finns ett område med byggnader, cirka 35 m långa och upp till 9 m brett, åtminstone fyra ruiner några meter ifrån varandra, tre av dem ligger tillsammans men den yttre ligger lite åtskild. 
Den sydligaste ruinen är otydlig vid väggränsen, men det är tydligt att det finns människoverk i marken." 
(Byggðasögu Skagafjarðar IV, Skagafjörðurs bygdehistoria volym 4, s. 172-173.) 
Ytterligare beskrivning: 
Den forntida gården Risamýri i trakten av Réttarholt i Akrahreppur. 
Sett mot sydost över den övervuxna Skiphóll.
Beskrivning:
Miðhúsaselland är det första fårbetet ii Deildardalursbygden, på västra sidan, det enda som inte ligger i Vesturdalur eller Austurdalur/Seljadalur. 
Det sträcker sig från Háleggstaðamerkjar till Bjarkará, mittemot Tungufjallssporður. 
Dess norra gräns anges i Miðhúss markgränsbrev. 
"Nedanför och utåt mot Háleggsstaðir, från skyddet vid kanten av Afréttará. 
Därifrån, raka vägen till Grænadragur och sedan så långt man kan se till passet på bergskanten utanför Bjarkarskálur." 
1709 slutade Miðhúsabændur att ha fäbod i Deildardalur. 
Fastighetsregistret säger: "Fäbod i Deildardalur i väster där marken kallas Björk, men kan inte användas för att den ligger för långt bort förutom för de mäktiga männen." 
Miðhúasel ligger cirka 405 meter utanför Bjarkará, på en lång ås nere på slätten vid foten av sluttningen, mittemot gården i Stafn. 
Söder om kullen finns ganska tydliga fäbodsruiner och en kort bit därifrån finns 8 meter långa fårfållor. 
Norr om kullarna finns andra fäbodsruiner, tre stycken, totalt cirka 16 meter långa. 
(Byggðasögu Skagafjarðar VII, Skagafjörðurs bygdehistoria volym 3, Hofshreppur, 186).  
Ytterligare beskrivning: 
Översiktbild av ruiner vid Miðhúsasel. 
Sett söderut.
Beskrivning: 
Sedan 2003 har Byggðasafn Skagfirðinga och Byggðasaga Skagafjarðar, Skagafjörðurs bygdemuseum och bygdehistoria, ansvarat för ett gemensamt forskningsprojekt som syftar till att dokumentera och undersöka de äldsta resterna av Skagafjörður, med särskild tonvikt på trakten och traktens fjällområden. 
Från början har projektet varit en del av arbetet med att skriva Byggðasagan, Byggdehistoren, nu har fyra framgångsrika volymer publicerats. 
Byggðasagan skiljer sig från andra lokalhistoriska böcker genom att det läggs större vikt vid gårdarnas forntida historia och studiet av alla typer av arkeologiska lämningar som kan läggas till deras historia. 
De två sista volymerna av Byggðasagan innehåller detaljerade kapitel om forntida bosättningar i de inre dalarna i Austurdalur och Vesturdalur, där historien är sammanflätad med resultaten av arkeologiska utgrävningar som har ägt rum på utvalda platser. 
Resterna av en gammal bondgård, den så kallade Gerði (65°35'315/19°18'940), ligger cirka 400 meter ovanför byn i Flugumýrarhvammur. 
Det har länge legat ett [avskilt beläget] fårhus där och gjorde så fram till 1960-talet. 
1856 fanns det 30 fårhus i gott skick. 
Ett litet tun var inhägnat och slogs där fram till mitten av 1900-talet. 
Ruiner av två [avskilt belägna] fårhus kan ses, men tydligt synliga lämningar av mänskliga boningar finns i ett betydligt större område än runt fårhuset. 
Senast stod här dock bara ett fårhus, det som syns i den södra ruinen. 
Det har bildats en betydande gräsmarksbank och det syns en liten kulle i backen, men en mycket hög höjd blockerar utsikten mot norr. 
Här är gårdsnamnet Hvammur naturligt eftersom området bildar en bred dal. 
Sluttningen nedanför kallas Hallið men man ser inte från gården och upp i dalen. 
Upp från Gerði, högre upp i backen, finns det några framträdande sandkanter och klippblock och vatten rinner ner i en bäck som här kallas Gerðisklauf. 
Den rinner norr om Gerði och är även gårdsvatten till hemmanet i Flugumýrarhvammur. 
En större forntida gärdesgård finns i söder, över och ner norrut litegrann, den verkar gå en bit bortom bäcken så att brunnen skulle kunna ligga inom gärdesgården. 
Bäcken går cirka 40 meter utanför den antagna gårdskullen. 
Längst ner är det inte möjligt att med säkerhet skilja gärdesgården från myrmarken nedanför. 
Det finns ruiner på tre ställen. 
Först och främst lämningar efter ett [avskilt beläget] fårhus som utan tvekan har byggts ovanför gården, eftersom detta är den bästa platsen för ett hus och bildar en liten gårdskulle (65°35'315/19°18'940) med rester av byggnationer över ett större område. 
Forntida ruiner ligger direkt söderut, söder om gärdesgården (65°35'300/19°18'915). 
Längst ner på tunet, på en liten kulle nedanför gårdskullen, ligger det tredje ruinområdet (65°35'296/19°18'958). 
Det fanns ett baggehus ordagrant vid de [avskilt belägna] fårhusen på 1900-talet, men ruinerna där är mycket större än motsvarigheten till ett baggehus. 
Det är våtmark framför kullen och gärdesgården har troligen legat under den. 
Bosättningen i Gerði har för länge sedan fallit i glömska och därmed även gårdens namn. 
Fastighetsregistret från 1713 berättar om denna plats: "Fårhusplatsen är omgiven som om det en gång varit bebyggt där. Ingen vet något mer om det." 
(Árn Magnússons och Pál Vídalíns Jordabok IX, s. 187). 
Det finns olika tecken på att det här är den äldsta platsen för gården, gården Hvamm, som sedan dess har flyttats därifrån och ner ut ur dalen, men namnet blev kvar (Byggðasögu Skagafjarðar IV, Skagafjörðurs bygdehistoria volym 4, s. 145-46). 
Ytterligare beskrivning: 
Översikt över Gerður, en gammal gård i Flugumýrahvammur i Akrahreppur. 
Sett västerut. 
Héraðsvötn kan ses högst upp på bilden och gården längst till höger är Réttarholt. 
Beskrivning: 
Spáná är den innersta gården i Unadalur, norr om Unadalsá. 
Där finns betydande gårdsruiner, fortfarande mycket tydliga, och en hel del uthusruiner över hela fältet och bortom det. 
Vallmuren är kraftig ovanför ängen under Spánárhóll, den främre delen är belagd med torv och den yttre delen är gjord av sten och når cirka hundra meter ner till skredgrunden. 
Tunet har varit ganska stort, på torr torvmark och övervuxna jordskredslager i Spáná, hård mark som är svår att bryta. 
Spáná övergavs 1921 och det finns inte längre några hus kvar. 
Marken ägs nu av Upprekstrarfélag Unadalsafréttur, Unadalurs fjällbetessamfällighet och är en del av Unadalurs betesmarker (Veðmálaskrár, Inteckningsregistret, nr. 4756). 
Spáná verkar ha legat öde under lång tid under medeltiden. 
Det är okänt när området först bebyggdes, men biskopssätet i Hólar verkar ha förvärvat marken på 1400-talet. 
Marken är tidigast dokumenterad i biskopssätets register från 1525 och räknas där som obebyggd ödemark (Diplomatarium Islandicum, Íslenskt fornbréfasafn, 302). 
Källan hävdar att Þorbergur Bessason, häradshövding på Hof, hyrde Spáná från Hólar i mitten av 1500-talet och hade en fäbod där medan han drev gården på Hof (Jarðabréf á Þjóðskjalasafni, Markhandling i Islands Nationalarkiv, 2 (72) B). 
Marken har byggts upp igen under andra hälften av 1600-talet, eftersom den omnämns i biskopssätet i Hólars förteckning 1666 och i Jordaboken 1709 står att den byggdes upp från ödemark för 40 år sedan, d.v.s. någon gång före 1670 (Árn Magnússons och Pál Vídalíns Jordabok, 247). 
I Jordaboken 1709 uppskattas Spáná bara till 6 hundraden och det är ett lågt mått som utan tvekan beror på markträngsel och stor osäkerhet. 
I Johnsens Jordabok från 1847 sägs marken vara 6 hundraden, men fotnoten från distriktskommissionären värderas den till 8 hundraden (Árn Magnússons och Pál Vídalíns Jordabok, 247; Johnsens Jordabok 1847, s. 270). 
År 1849 var "Spáná bondeegendom i nuläget 8 hundraden" (Jordabok 1849 nr. 78). 
ommaren 2013 togs ett antal borrkärneprov i Spáná. 
Det fanns spår av en bosättning redan på 1000-talet, kanske tidigare. 
Bosättningen kan ha övergivits redan på 1100-talet. 
Det kan dock ha varit en viss byggnation där, kanske var det fortsättningsvis en fäbod efter det att bosättningen upphörde på 1100-talet och innan den byggdes upp igen på 1600-talet.  
Ytterligare beskrivning: 
Kári Gunnarsson i en stugruin öster om fårhusruinen. 
Sett mot nordost. 
Beskrivning: 
Hrappsá var ett arrende till Skuggabjarg och stod norr om floden med samma namn i Deildardalur i väster, mellan Skuggabjarg och Stafshóll. 
Det är osäkert hur stor mark arrendatorn hade, annat än tunet, som avgränsas av en gammal gärdesgård. 
Olyckligtvis finns inga kvarvarande skriftliga källor om Hrappsás existens före 1831, förutom en folklegend som verkar ha sitt ursprung i de första århundradena av de isländska bosättningarna. 
Dessa legender hittades i handskrifter från åren 1368 och 1428, som tyvärr gått förlorade (HSk. 403. fol. Platsnamnbeskrivning från Deildardalur. Jón H. Árnason). 
Hrappsá nämns inte i fastighetsregistret 1709, vilket måste betraktas som ganska ovanligt, men kan ha sin förklaring (Árn Magnússons och Pál Vídalíns Jordabok X, s. 209-210). 
Skuggabjörg var öde 1709 och därför fanns ingen boende i området som kunde rapportera om de lokala förhållandena. 
Hrappsá verkar ha glömts bort. 
Ólafur Olavius reseskildring från 1777 nämner inte heller Hrappsá i listan över ödegårdar i Hofshreppur.  
Gården var bebyggd från 1831 och beboddes till och från fram till 1872, då Hrappsá övergavs och har inte varit bebodd sedan dess. 
Hrappsá nämns i en fotnot i Johnsens förteckning över gårdar från 1847, där det står att prästen nämner arrendet Hrappsá, men närmare information om gården finns inte och därför finns den inte med i själva förteckningen (Jarðatal Johnsen, Johnsens förteckning över gårdar, 1847, s. 270). 
Platsen för gården ligger nära och ovanför vägen (västra Deildardalsvegur) som går mellan Skuggabjargar och Stafshóll, direkt framför Hrappsárskrið. 
Tunet ligger i en liten sluttning, välväxt och tjock och har aldrig jämnats ut. 
Innanför gärdesgården finns några tydliga ruiner från en bostad på 1800-talet men även grunder för äldre ruiner. 
Färdvägen till Hrafnsá har legat långt från gården när den första gården byggdes och idag har en del av tunet och gärdesgården hamnat under flodskred. 
Det går inte att säga när skredet gick över tunet och förstörde gärdesgården. 
Det är dock uppenbart att invånarna i Hrappsá på 1800-talet inte har haft någon anledning att återställa den. 
Gården har uppenbarligen tagit sitt namn från floden som ligger bredvid, den har länge kallats Hrappsá men har under senare år ändrats till Hrafnsá. 
I ortnamnsregistret från 1938 används namnet Hrappsá, men i mark- och personregistret, Jarði og búendatal, från 1953 heter gården Hrafnsá. 
I församlingsbeskrivningen från 1839 anges att bredvid Hrappsá står den nya gården Hrappsá (Läns- och församlingsbeskrivningar, Sýslu og sóknarlýsingar II, s. 137).  
Under 1900-talet kallades Hrappsá för Hrafnsárkot. 
Ortsnamnsregistret anger att namnet Hrafnsárkota används av lokalbefolkningen i dagligt tal (Rósmundur Ingvarssons ortsnamnslista, Örnefnaskrá Rósmundar Ingvarssonar). 
Profil 1. 
En profil togs fram i den norra delen av gärdesgården, där en bulldozerväg hade bildat ett perforerat snitt i den. 
Profilen rensades och grävdes upp cirka 40 cm nedanför gården för att komma ner i orörda jordlager.
 Profilen visade en 50 cm hög torvvägg som har byggts efter 1104. 
H1104-pyroklastern verkade orörd under väggen, men under fanns torv rotad med H3-pyroklastern, cirka 8-10 cm tjock hög. 
Det är vanligt att torv och jord används för att täta under väggar så att underlaget blir så jämnt som möjligt, vilket kan förklara gräsrötterna. 
Å andra sidan måste det anses vara ganska intressant att vulkanen 1104 tycktes ligga orörd över den. 
Så askan har fallit under den tid då muren byggdes. 
Det är dock inte uteslutet att skiktet låg längst ner i den torv som användes för att täcka det tvärgående hålet som grävdes. 
Det är dock klart att gärdesgården iordningställdes först efter pyroklaster-nedfallet 1104, men profilen visade inte avgörande tecken på annan pyroklaster, vare sig i gräset eller ovanför gården. 
Profil 2 
En annan uppblåst profil togs fram i den yttre delen av gärdesgården. 
Där fanns jordlager som liknade dem i profil 1, förutom att marken uppenbarligen hade iordningställts efter år 1300. 
Pyroklaster från Hekla-1300 fanns i den översta torven i marken. 
Det var inte möjligt att bestämma jordlagret längst ner på väggen, eftersom vatten ackumulerats längst ner i profilen, då en bäck från myren utanför gården här rann genom väggen. 
Tolkning: 
Det är tydligt att den första bosättningen på Hrappsá är från 1000-talet, kanske tidigare, och där en stuga, fårfålla och halvcirkelformat markskikt är de äldsta lämningarna inom tunet. 
Gärdesgården indikerar dock att Hrappsá var bebott efter 1104, kanske ända fram till 1300-talet. 
Lämningar från den bosättningen ligger antagligen under resterna av 1800-talets bosättning. 
Det är dock tydligt att gården har varit öde under lång tid innan den byggdes om under några decennier på 1800-talet. 
Ytterligare beskrivning: 
Markprofil från norra delen av gärdesgården på Hrappsá. 
Sett uppifrån. 
Beskrivning: 
Marken för de lägsta fårmarkerna i den västra delen av Unadalur tillhörde Þönglaskáli på Höfðastrand. 
Den mäter ca. 180 hektar. 
Gränsen för Þönglaskálaselland i norr, mot Bjarnastaðagarður, är enligt en markgränsbok från år 1890, "vid Puntskriða, på väg uppför fjället." 
Jóhann Ólafssons ortnamnsregister innehåller en mer detaljerad beskrivning av dessa gränser: "Från markgränsen till Bjarnastaðagarður, som utgjordes av stor sten vid Unadalsá, vid stranden av den så kallade Puntskriða, rakt mot Kisukinn nedanför fjällstugan Kisa och rakt upp på fjället." 
Þönglaskálasel ligger väster om Unadalsá, på en mycket hög bank, mittemot Spánás fårfållor. 
Det finns rester av byggnader på minst sju platser, några mycket gamla, andra tydligt mycket yngre. 
Huvudruinen liknar inget annat än en gårdsruin. 
Det finns i sju avdelningar och vegetationen i den är mycket kraftigare och grönare än omgivningens, vilket indikerar att den inte kan vara mycket äldre än 200 år, högst 300 år. 
Cirka 12 meter ovanför finns ruiner av små fårhus. 
På fyra andra platser finns ruiner av småhus eller fårfållor (...). 
Sommaren 2013 genomfördes en mindre arkeologisk utgrävning med en kärnborr vid Þönglaskálasel. 
Det visade sig vara svårt att få tillfredsställande resultat eftersom borren ofta fastnade i sten innan den nådde ner till en acceptabel nivå. 
Det var därför inte möjligt att bestämma åldern på gårdsruinen. 
Men dess skick och askan från 1766 indikerar att väggarna byggdes om efter 1766 års utbrott. Under dessa husruiner visade det sig dock finnas en annan byggnad, kanske lämningarna av en fäbod eller ett gårdshus. 
Vid sidan om fanns otydliga och nersjunkna väggar från äldre byggnader där det var möjligt att identifiera åtminstone två utrymmen. 
Det visade sig vara byggnaden av ett hus som antagligen hade rivits 100-200 år innan gårdshuset byggdes ovanpå och vid sidan om. 
Ett tätt, moaskerikt golv med en kolrester som tydligt har varit i en människobostad. 
Cirka 15 cm orörd lössjord låg ovanpå dessa lämningar. 
Torven som visade sig i kärnprovet innehöll pyroklaster från Heklas utbrott 1104 och väggarna har byggts efter utbrottet. 
Det är möjligt att utläsa lämningar från tre bosättningsperioder där. 
En arkeologs tolkning var att det ursprungligen fanns en fäbod, byggd efter 1104 men troligen övergiven på 1300- eller 1400-talet. 
Ruiner av en stuga kan vara knutna till en fäbod eller boskap på platsen efter det att den äldre fäboden övergivits. 
På 1700- eller 1800-talet fanns där en kortlivad bosättning. 
En lokalhistoriker minns att han hört någon prata om Þönglaskálagarður. 
Det kan ha varit namnet på gården som låg där under en kort tid på 1700-talet eller i början av 1800-talet, men inga registrerade källor har hittats. 
Det är i varje fall inte en beboelig plats när vad gäller tillgång på ängar och gräsmarker, men fäbodsplatsen är beboelig. 
(Skagafjörðurs bygdehistoria - Byggðasaga Skagafjarðar VII. Hofshreppur, 268). 
Ytterligare beskrivning: 
Uthusruiner ovanför gårdshusruinerna vid Þönglaskálasel. 
Sett mot nordost.
Beskrivning: 
Ödebygd och dalar III. 2008. 
Hólakot i Viðvíkur i Viðvíkur-trakten. 
Hólakot omnämns tidigast i källor tillsammans med Viðvík och Kvígildis¬hóll i förvaltningsberättelsen för biskopssätet i Hólar från 1388 där mark som ägs av biskopssätet är listad (Diplomatarium Islandicum, Íslenskt fornbréfasafn, III: 410). 
I en annan lista över Hólastaðurs ägor från 1449 listas Viðvík tillsammans med Hólakot (Diplomatarium Islandicum, Íslenskt fornbréfasafn, V: 36, 43). 
I Margeir Jónssons ortsnamnsregister står i sista stycket: "Hólakot, som är en forngammal gård - ligger i Viðvíkurland men byggdes om 1920. 
Den forntida värderingen av Hólakot var 20 hundraden. och omkring år 1388 var hyran. 3 tre märken vadmal. 
Genom kungligt dekret den 8:e maj 1805 placerades Viðvík "tillsammans med stugan" som en bostad för distriktskommissionären och den har följt med huvudmarken ända sedan dess. "
(Viðvíkurs ortnamnregister - Örnefnaskrá Viðvíkur Margeir Jonsson registrerade. Isländska ortsnamnsinstitutet - Örnefnastofnun Íslands s. 3). 
Sverrir Björnssons ortnamnsregister säger: "Ovanför sundet [Hólakotssund] finns en liten stuga som heter Hólakot, med hänvisning till Margeir Jónssons beskrivning 
(Viðvíkurs ortnamnregister - Örnefnaskrá Viðvíkur Sverrir Björnsson registrerade. Isländska ortsnamnsinstitutet - Örnefnastofnun Íslands s. 3). 
Hólakot kan ha varit bebodd 1921-1934. 
I Hólakot kan du se resterna av en gärdesgård och byggnadsresterna från de båda stugor som stod där senast, men det finns även stora fornlämningar på gärdesgården som det inte finns några källor till. 
Totalt tre marksnitt gjordes vid Hólakot, förutom att ett antal kärnprover togs för vidare analys av lämningarna.  
Ytterligare beskrivning: 
Hólakot marksnitt 2. 
Den forntida gården Hólakot i Hjaltadalur. 
Marksnitt 2 togs i gärdesgårdens norra del. 
Det hittades minst två byggnationsperioder på gården. 
Det verkar som att gården delvis kollapsade när pyroklastern från vulkanutbrottet 1104 nedföll. 
Det är möjligt att gården byggdes upp igen, men inga pyroklaster hittades ovanpå själva gården och det fanns inga tecken på 1104-pyroklaster i torven. 
Den nedre delen av gården var byggd av torv som innehöll fint svart pyroklaster- det kan vara ett pyroklasterlager från Vatnajökull som nedföll omkring 1000 e.Kr.
Beskrivning: 
Bjarnastaðir är en ödegård på östra sidan av Unadalur, 140 meter över havet. 
Marken ligger mellan Bjarnastaðaá och utsidan av Tungufjall och Spánárdalur och Spáná framför. 
Runt marken ligger Grundarland utanför, högt fjäll ovanför, Spáná på insidan och Unadalsá nedanför mittemot Þönglaskálaselland och Bjarnastaðagarður. 
Bjarnastaðir omnämns tidigast i källor 1449, då marken ägdes av biskopssätet Hólar. 
Gården ödelades 1947 och alla hus där har för länge sedan förfallit. 
Marken avsattes formellt till betesmark 1961 (Skagafjörðurs bygdehistoria volym 7, Byggðasaga Skagafjarðar VII, 281).    
Ytterligare beskrivning: 
Gärdesgården vid Bjarnastaðir. 
Sett mot nordväst. 
Beskrivning: 
Hagakot är en ödegård och det var den främsta gården i Hjaltadalur öster om floden under de senare århundradena. 
Marken var inte en självständig gård på 1800-talet, utan en slags bondgård under Hólar och den hade inga specifika gränser. 
Den var bebodd 1862-1888. 
Gården stod i den norra änden av Hagafjall, direkt nedanför Tröllkonusætur, som är ett klippsediment längs den mellersta sluttningen norr om bergskedjan. 
Vid Hagakot finns det tre ruiner av [avskilt belägna] fårhus och det finns fortfarande ett fårhus kvar som byggdes i mitten av 1900-talet. 
Längst bort och nederst på det gamla tunet finns en ruin som inte verkar ha varit ett nyttohus. 
Ruinen var uppdelad i fyra delar och borrkärneprov togs i dess väggar och golv.
Tolkning av kärnprovet: Spår av en eldstad indikerar att detta varit en människobostad. 
Den var troligen bebodd på 1600-talet, möjligen fram till 1700-talet. 
Ytterligare beskrivning: 
Rester av ett boningshus vid Hagakot i Hólahagi. 
Sett från nordväst.
Beskrivning: 
Bäcken omnämns först i mitten av 1300-talet, men arkeologiska fynd indikerar att området var bebott från de tidigaste bosättningstiderna. 
Jordbruket upphörde 1958 och marken är nu en del av Ennis mark och nyttjas därifrån (Byggðasaga Skagafjarðar V, Skagafjörðurs bygdehistoria Volym 5, s. 269-270). 
Inga fler byggnader är uppförda, men gårdskullen är fortfarande tydligt igenkännlig. 
Gärdesgården kan ses delvis till väster och norr om gårdskullen och det finns två ruiner vid dess västra del. 
Cirka 20-50 meter direkt norr om gårdskullen finns otydliga fornlämningar, ruiner av stugor och andra byggnadsrester. 
Borrkärneprov togs i ruiner och gärdesgård, förutom att ett marksnitt togs inne i stugruinerna. 
Ytterligare beskrivning: 
Lækur i Viðvíkursveit. 
Marksnitt 1 i stugruin, botten på marksnittet. 
Ett marksnitt togs i den östra delen av ytterväggen av ett långsträckt bostadshus eller stuga söder om Lækjars eget gårdstun. 
Cirka 5 cm under gräsrötterna [1] fanns orörd pyroklaster H1300 men ingen människobostad kunde ses i lössjorden [2] ovanför den. 
Mellan 1300 och 1104, som också det var orört i profilen, fanns det ett lager lössjord [3] med några spår av 1104 och en spridd moaska, men annars mycket små tecken på en människobostad. 
H1104 låg i cirka 2 cm tjocka skikt ovanpå en torvvägg som skönjdes till väster om diket och var något mer otydlig längs hela profilen. 
Cirka 2 cm orörd lössjord [4] fanns mellan pyroklastern och den övre delen av torvväggen, med ett upp till 20 cm tjockt lössjordskikt [4] över en kollaps av väggen [5] men den har rasat åt öster  
Byggnaden verkar därför ha övergivits strax före 1104 års vulkanutbrott, men det är inte möjligt att ange med större noggrannhet när den byggdes. 
Tolkning: 
Byggnaden övergavs något tidigare än 1104, och dess murar verkar då ha kollapsat. 
Borrkärneproven indikerade att det varit ett bostadshus och formen på ruinen indikerar också att det var en stugruin. 
Det finns få bevis på människobostad efter det att huset kollapsade eller jämnades under 1104 års vulkanutbrott. 
Det är osäkert om detta innebär att det funnits en bosättning där, men åtminstone verkar gårdstunet inte ha legat på samma plats. 
Det finns ytterligare bevis för bosättning mellan 1104 och 1300, men inte överväldigande många. 
Beskrivning: 
År 2013 undersöktes ett antal platser i den forntida Hofshreppur i samband med projektet "Öde bosättningar och dalar i Skagafjörður", Eyðibyggð og afdalir Skagafjarðar (VII). 
Tyngdpunkten lades på lämningar i Deildardalur och Unadalur och huvudsyftena var följande: 
att söka efter och lokalisera forntida gårdar, fähus och andra lämningar som kan ge kunskap om landsbygdshistorien i Skagafjörður. 
att undersöka åldern på utvalda lämningar med marksnitt och/eller borrkärneprov tagna i marken och ruinernas ytterväggar för att bestämma ålder och eventuellt byggnadsstadium. 
Kärnprover togs även från golven för att avgöra om det varit människobostäder. 
Att presentera och uppmärksamma lämningarna så att de kan beaktas vid planering och konstruktion. 
Ytterligare beskrivning: 
Sett in i Unadalur från Svínavellir. 
Sett österut.
Beskrivning: 
Hrappsá var ett arrende till Skuggabjarg och stod norr om floden med samma namn i Deildardalur i väster, mellan Skuggabjarg och Stafshóll. 
Det är osäkert hur stor mark arrendatorn hade, annat än tunet, som avgränsas av en gammal gärdesgård. 
Olyckligtvis finns inga kvarvarande skriftliga källor om Hrappsás existens före 1831, förutom en folklegend som verkar ha sitt ursprung i de första århundradena av de isländska bosättningarna. 
Dessa legender hittades i handskrifter från åren 1368 och 1428, som tyvärr gått förlorade (HSk. 403. fol. Platsnamnbeskrivning från Deildardalur. Jón H. Árnason). 
Hrappsá nämns inte i fastighetsregistret 1709, vilket måste betraktas som ganska ovanligt, men kan ha sin förklaring (Árn Magnússons och Pál Vídalíns Jordabok X, s. 209-210). 
Skuggabjörg var öde 1709 och därför fanns ingen boende i området som kunde rapportera om de lokala förhållandena. 
Hrappsá verkar ha glömts bort. 
Ólafur Olavius reseskildring från 1777 nämner inte heller Hrappsá i listan över ödegårdar i Hofshreppur.  
Gården var bebyggd från 1831 och beboddes till och från fram till 1872, då Hrappsá övergavs och har inte varit bebodd sedan dess. 
Hrappsá nämns i en fotnot i Johnsens förteckning över gårdar från 1847, där det står att prästen nämner arrendet Hrappsá, men närmare information om gården finns inte och därför finns den inte med i själva förteckningen (Jarðatal Johnsen, Johnsens förteckning över gårdar, 1847, s. 270). 
Platsen för gården ligger nära och ovanför vägen (västra Deildardalsvegur) som går mellan Skuggabjargar och Stafshóll, direkt framför Hrappsárskrið. 
Tunet ligger i en liten sluttning, välväxt och tjock och har aldrig jämnats ut. 
Innanför gärdesgården finns några tydliga ruiner från en bostad på 1800-talet men även grunder för äldre ruiner. 
Färdvägen till Hrafnsá har legat långt från gården när den första gården byggdes och idag har en del av tunet och gärdesgården hamnat under flodskred. 
Det går inte att säga när skredet gick över tunet och förstörde gärdesgården. 
Det är dock uppenbart att invånarna i Hrappsá på 1800-talet inte har haft någon anledning att återställa den. 
Gården har uppenbarligen tagit sitt namn från floden som ligger bredvid, den har länge kallats Hrappsá men har under senare år ändrats till Hrafnsá. 
I ortnamnsregistret från 1938 används namnet Hrappsá, men i mark- och personregistret, Jarði og búendatal, från 1953 heter gården Hrafnsá. 
I församlingsbeskrivningen från 1839 anges att bredvid Hrappsá står den nya gården Hrappsá (Läns- och församlingsbeskrivningar, Sýslu og sóknarlýsingar II, s. 137).  
Under 1900-talet kallades Hrappsá för Hrafnsárkot. 
Ortsnamnsregistret anger att namnet Hrafnsárkota används av lokalbefolkningen i dagligt tal (Rósmundur Ingvarssons ortsnamnslista, Örnefnaskrá Rósmundar Ingvarssonar).  
Ytterligare beskrivning: 
Forntida fårfålla på Hrappsá. 
Sett norrut. 
Beskrivning: 
En arkeologisk undersökning utfördes på ett av arrendena till kyrkomarken Miklabær i Akrahreppur. 
Gårdens namn är okänt men denna diskussion finns i Byggðasögu Skagafjarðar IV, Skagafjörðurs bygdehistoria volym 4, där mark i Akrahreppur diskuteras. 
En av Miklabærs fyra gårdar var gården Jaðar. 
Fastighetsregistret 1713 nämner följande: "tredje arrendet, öde på samma sätt som det sägs om Miklabæjarkot..." 
År 1753-1757 bodde Jaður Grímur Jónsson och Guðrún Gottskálksdóttir från Hreiðarsstaðir i Svarfaðardalur, men hon var helsyster till Þorvaldur Gottskálksson, präst i Miklabær 1747-1762 och halvsyster till Gottskálk Blander i Mið-Grund. 
Namn på andra invånare i Jaðar är inte kända och det verkar som om prästen Þorvaldur har tillåtit sin syster och svåger bo och bygga på en gammal ödestuga (Svarfdælingar II, s. 96). 
Även om det låter konstigt så har nutida människor glömt var Jaðar arrende låg, eftersom de inte längre ser några direkta spår av det. 
Om man tittar på miljön måste en viss plats dock anses vara ganska sannolik utan att det finns riktiga några bevis. 
I det nordöstra hörnet av det gamla tunet som kallas Húsahóll, söder om Bæjarlækur och ovanför huvudvägen. 
Där böjer sig den gamla gärdesgården över kullen mot toppen. 
Där fanns ett fårhus fram till andra hälften av 1900-talet och det finns fortfarande tydliga tecken på två [avskilt belägna] fårhus som vetter utåt och söderut, sida vid sida med en lada mittemellan (65°30'500/19°17'575). 
Detta är i utkanten av tunet och en mycket trolig gårdsplats, med nära till bäcken. 
Men lämningar från forngårdar har hittats längst ner i Miklabæjarnes. 
Héraðsvatn har sedermera eroderat bort en del av tunet, kanske så mycket som upp till hälften av det. 
Det som återstår är en halvcirkel av den forntida gärdesgården och en liten del av gårdskullen. 
Det finns ett mycket gammalt ruinlager på ett ställe på gärdesgården, i nordost. Kanske är det en gammal stuga. 
En långsträckt kulle som Vötnin till största delen har eroderat bort och som är markerad B på bifogad ritning är grönare än omgivningen. 
Det ger en indikation på att en människobostad där inte är många århundraden gammal. Kanske är detta en gammal gårdskulle. 
Odlingar i sådana människobosättningar eller ruiner kvarstår i minst 200-300 år. 
Det är osäkert om den forntida gården är densamma som Jaðar som omnämns i Jordaboken eller om den handlar om en femte gård. 
Den 10:e juli 2007 genomfördes arkeologiska utgrävningar på platsen för åldersbestämning.. "(Hjalti Pálsson (red.) 2007: Skagafjörðurs bygdehistoria volym 4, Byggðasaga Skagafjarðar IV.   Akrahreppur. 
Sögufélag Skagfirðinga - Skagfjörðurs historiska sällskap Sauðárkrókur). 
Ytterligare beskrivning: 
En namnlös gammal gård på Miklabærs mark i Akrahreppur. 
Två marksnitt togs, den ena i gärdesgården och den andra i en ruin. 
Gärdesgårdsmuren är lagd efter år 1300, men det fanns ingen pyroklaster ovanför den, så det var inte möjligt att fastställa den övre åldersgränsen. 
Detsamma kan sägas om ruinen där ett marksnitt gjordes, det var inte möjligt att avgöra om det byggdes där före år 1300. 
Gården var därför troligtvis bebodd efter 1300 men var öde innan Árn Magnússons och Pál Vídalíns Jordabok skrevs 1713.
Beskrivning: 
Kärnproverna togs i ruinerna av Grafarsel i Deildardalur. 
Det finns betydande lämningar från fårhuset, både av äldre fårhus och resterna av en gård som fanns där i mitten av 1800-talet. 
Grafarsel ligger cirka 450 meter innanför Bjarkará, nere vid stranden av Grafará.  
Seljadalur nämns tidigast i en köpehandling från slutet av 1300-talet och namnet är utan tvekan gammalt. 
Det är inte osannolikt att bönder nere i dalen eller på Höfðastrand redan under de första bebodda århundradena hade fårhus runt bosättningen i Deildardalur (Diplomatarium Islandicum, Íslenskt fornbréfasafn III, s. 488). 
Pastor Páll Erlendsson säger om fårhus i Deildardalur i en församlingsbeskrivning från 1839: "All Óslandshlíðs mark, Gröf, Enni och Hof [har [avlägset belägna] fårhus], de två sista i Unudalur, de andra i Deildardalur. 
Inget av dem används nu, utom av Gröf, en månad varje sommar. 
De har övergivits på grund av avståndet, många relaterade svårigheter och har hittills aldrig varit lönsamma. 
Människor gräver efter kol där och driver kastrerade får och otämjda hästar dit, och jordbruksmarken är inget annat än själva fårhusmarken [...] "(Sýslu- og sóknalýsingar Skagafjarðarsýslu, Skagafjörður härads läns- och sockenbeskrivning, s. 139). 
De tydligaste lämningarna är resterna av en gård från 1800-talet som delvis ligger ovanpå resterna av äldre byggnader. 
Ruinerna av den yngsta gården ligger överst av lämningarna på en liten kulle och det fanns spår av tre utrymmen i gården, men de mest etablerade öster om gården var resterna av en grönsaksträdgård. 
Ruinerna av en hydda ligger några meter söder om grönsaksträdgården och härrör från den senaste användningsperioden. 
I ruinerna som gården står på kan du se åtminstone tre fack. 
Strax öster om den fanns en slags nedgrävning. 
Cirka 8 meter nordost om grönsaksträdgården fanns resterna av ett äldre fårhus, men inga yngre byggnader fanns ovanpå den. 
I den fanns åtminstone tre utrymmen och bifogade fårfållor. 
Ruinerna stod mycket nära kanten ovanför floden och var därför utsatta för erosion. 
Väggarna var väl nedsjunkna i jorden. 
Flera kärnprov togs i lämningarna. 
De flesta slog direkt i sten under ytan, eftersom det fanns många stenar i väggarna i både yngre och äldre ruiner. 
Det var inte möjligt att bestämma åldern på lämningarna i de tre kärnproverna som man lyckades ta där. 
Cirka 4 meter norr om fårhusruinen fanns långsträckta fårfållor som tillhörde fårhusruinen. 
Cirka 30 meter direkt norr om den yngsta gårdsruinen fanns resterna av två uthus, ett fårhus och en ladugård. 
De förstörda murarna i uthusen var i gott skick och det var uppenbart att det funnits en gård vid fårhusen. 
Dessa uthus var från 1800-talets gård. 
Tolkning. 
Det var inte möjligt att uppskatta åldern på lämningarna i Grafarsel. 
Ytterligare beskrivning: 
Sett ut över ruinerna i Grafarsel. 
Sett österut.
Beskrivning: 
En otydlig gård som går från öster till väster över Ástunga mellan Kolbeinsdalsá och Hjaltadalsá i Skagafjörður.  
Ytterligare beskrivning: 
Gårdsskikt mellan Hjaltadalsá och Kolbeinsdalsá i Skagafjörður. 
Sett från nordost. 
Beskrivning: 
I Ólavíus reseskildring (Ólafur Olavius (1965)) omnämns gården Ytri-Heljará och det står att den förstördes av en översvämning. 
Heljarár omnämns även i Gudmundur den Godes saga. 
Gårdens läge har varit okänt, men under forskning i samband med skrivandet av Byggðasagan undersöktes fäbodar i trakten av Bjarnastaðir, vid floden Heljará. 
Ytterligare fältforskning sommaren 2008 avslöjade, förutom uppenbara fäbodsruiner, resterna av äldre lämningar. 
Ruinerna ligger i den norra delen av flodselet, men det är tydligt att Heljará tidigare har runnit norr om selet, men rinner nu söder om det. 
Vid närmare granskning visade det sig att floden har svept bort några av de äldre ruinerna, det var dock möjligt att dämma upp en profil i flodbanken för att ytterligare undersöka lämningarna. 
Ytterligare beskrivning: 
Lämningar vid stranden av floden Heljará i Kolbeinsdalur. 
Sett mot sydost.
Beskrivning: 
Stafshóll ligger vid mynningen av Deildardalur i söder men ansågs antagligen höra till Höfðastrandur. 
Stafshóll sägs nu allmänt vara den lägsta gården i Deildardalur, söder om Deildardalsá. 
Gården står i nordväst i den så kallade Stafshólsöxl. 
Gårdens namn skrivs antingen Stafshóll eller Stafnshóll. 
De äldsta källorna om gården finns troligen i Landnamsboken, som berättar historien om Oddleif. 
Hans föräldrar var Hrafna-Flóki och Gró, hans syster Höfði-Þórðar, men Oddleifur bodde på Stafshóll och delade den med Hjaltason på Hof i Hjaltadalur. 
Landnamsboken nämner även Arnór, son till Nafar-Helgi, en bosättare vid Grindli i Fljóti, Arnór slogs med Friðleif på Stafshóll. 
Stafshóll är därför utan tvekan det ursprungliga gårdsnamnet (Islänningasagorna del 1, s. 151). 
Marken har utan tvekan varit privatägd i många århundraden, men Oddleifur Stafur, Hrafna-Flókason, verkar ha varit den första ägaren enligt Landnamsboken. 
Namnet på marken finns inte i biskopssätet Hólars förvaltningsredogörelse från 1388 och förmodligen blev det inte biskopssätets egendom förrän på 1400-talet. 
Stafshóll var en av de marker som biskoparna i Hólar rådde över och ofta köpte och sålde. 
Marken ansågs tidigare århundraden vara värd 24 hundraden men på 1600-talet och senare värderades den till 20 hundraden (Árn Magnússons och Pál Vídalíns Jordabok IX, s. 239). 
I Jordaboken från år 1709 nämns ett arrende från Stafshóll, som redan då var öde: "Hjáleigugrey har varit här en gång och den enda höskörden som bonden på hemmanet tog hem, tror folk vara 20 eller 30 alnar. 
Inget kan byggas här igen utan att vara till nackdel för marken" (Árn Magnússons och Pál Vídalíns Jordabok, s. 239). 
Förmodligen har detta arrende varit det som kallats Stafshólsstekkur strax nedanför Stafshól. 
Det finns en tydlig gärdesgård runt två byggnadsskullar. 
Resterna av 
gärdesgården [1] är ganska tydlig, upp till en meter hög och cirka 2 meter bred. 
De omger ett tun som är cirka 100 meter långt från nordväst till söder och cirka 60 meter där det är som bredast. 
Ett otydligt gårdsområde [3] verkar korsa området strax söder om en möjlig gårdskulle. 
Om tunet någonsin har utökats eller minskats eller delats av bör vara osagt. 
Som nämnts tidigare finns det två kullar på tunet.  
Den västra kullen är en trolig gårdskulle, 21x6 m stor, men formar inte de tydliga konturerna av byggnader på den, men bulor i kullen indikerar att det har funnits en tvådelad eller tredelad ruin där [2].  
På den andra kullen söder om tunet finns två dubbla ruiner, troligen de högsträckta ruinerna som området har fått sitt namn från. 
Ruinerna ligger parallellt med den större i sydväst, cirka 11x3 meter stor. 
Fast nordost om det finns en mindre ruin 8x4m stor. 
Båda ruinerna är uppenbarligen mycket yngre byggnader än gärdesgården och ruinerna på den omnämnda gårdskullen.  
Strax väster om gärdesgården finns en otydlig gammal ruin 6x5 m stor och den är täckt med ljung. 
Kärnprover togs i en gärdesgårdsmur, en påstådd gårdskulle och en gammal ruin utanför gärdesgården. 
Endast fem borrkärneprov togs, eftersom resultaten var ganska enstämmiga. 
Gärdesgårdens kärnprov indikerade att den byggdes efter år 1104 men övergavs före år 1300 som låg orörd över gården. 
Detsamma gällde kärnprovet togs i gårdskullen, där resterna av människoboning, kol och moaska hittades. 
Ruinerna utanför gärdesgården verkar också ha kollapsat före år 1300. 
Vad gäller det "dåliga" arrendet som omnämns i Jordaboken hade det avskaffats ganska lång tid innan den skrevs. 
Det är dock inte uteslutet att det fanns vissa bosättningar där under en kort tid efter det att gården som gärdesgården tillhörde övergavs.  
Tolkning: 
Gården är avgränsad av en gärdesgård vid Stafshólsstekk har varit bebodd efter 1104 och gärdesgården har åtminstone kollapsat innan pyroklaster-nedfallet år 1300. 
Ytterligare beskrivning: 
Sett in i Deildardalur från Kotur i landet Stafn. 
Sett österut.
