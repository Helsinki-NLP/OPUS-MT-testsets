Denna uppsats är gjord på uppdrag av Tidningsutgivarnas organisation Tidningen i skolan och grundas på en kvantitativ enkätundersökning. 
Uppsatsen syftar till att försöka svara på den övergripande frågan "Vilka attityder har värmländska ungdomar till lokaltidningen?"
Enkäten ställde frågor om bakgrund, medievanor, och respondentens förväntningar på framtiden. 
Målgruppen avgränsades till gymnasieelever, och enkäten delades ut och samlades in under ett och samma besök i klasserna. 
De värmländska ungdomarna har generellt sett en relativt positiv bild av lokaltidningar. 
De allra flesta tror att de själva kommer att prenumerera någon gång i framtiden. 
Samtidigt visar resultaten att målgruppen spår lokaltidningarna en framtida nergång. 
Idag är det teven som är det främsta mediet för nyheter. 
Lokaltidningarna hamnar på en andraplats på samma lista. 
Får ungdomarna titta tio år in i framtiden tror de fortfarande att det är teven som är det främsta nyhetsmediet. 
Lokaltidningarna tappar på bekostnad av Internet, men hittas fortfarande på topp-tre.
Bara en tredjedel av ungdomarna upplever att deras lokaltidning riktar sig till deras åldersgrupp, knappt någon tvivlade på vuxna som målgrupp. 
När vi bad dem bedöma sina respektive lokaltidningars olika egenskaper var de flesta försiktigt positiva eller likgiltiga. 
Värmlands tidningar är enligt våra enkätsvar varken snygg eller ful, varken pålitlig eller opålitlig, och så vidare...
Resultatet ger en aning om att lokaltidningarna står inför, om inte sin död, så åtminstone en stor utmaning.
Syftet med detta arbete är att erhålla en ökad förståelse för på vilket sätt som relationsmarknadsföringssynsättet är närvarande i konsumentinriktade internetförsäljningsföretaget. 
En kvalitativ studie av fem företag inom konsumentinriktad internetvaruförsäljning genomfördes där företagens e-handelslösningar studerades och personal på företagen intervjuades. 
Resultatet visar att det i dessa företag verkar förekomma ett aktivt arbete med att etablera och underhålla relationer av främst monetär och social karaktär. 
Avseende relationsmarknadsföringssynsättet så förekommer begreppet, och synsättet finns till viss del etablerat bland några av de undersökta företagen.
Cochleaimplantat (CI) är en av de största medicinska innovationer som gjorts under de senaste 20 åren. 
Med hjälp av ett sådant kan barn med grav hörselnedsättning eller dövhet få möjlighet att höra och utveckla ett talat språk. 
Många barn med CI uppnår dock inte den förväntade språknivån. 
Orsakerna till detta är ännu inte fullt förstådda och vidare forskning är därför nödvändig. 
I föreliggande studie deltog 9 barn i åldrarna 6;7 – 12;4 år med CI. 
Syftet med denna studie var att undersöka kognitiv och språklig förmåga med fokus på arbetsminne och receptivt lexikon hos barn med CI. 
I detta syfte användes utvalda delar ur det datorbaserade testbatteriet SIPS (Sound Information Processing System) samt PPVT (Peabody Picture Vocabulary Test). 
Testresultaten analyserades på grupp- och individnivå. 
Dessutom jämfördes testresultaten med resultat från en kontrollgrupp normalhörande barn.
Barnen med CI presterade lägre än kontrollgruppen på gruppnivå. 
Enskilda individer presterade dock i nivå med barnen i kontrollgruppen vilket innebär att det är möjligt för barn med CI att uppnå goda resultat på de undersökta aspekterna. 
Resultaten i studien indikerar också att sen implantation inte alltid behöver vara ett hinder för god språklig utveckling. 
Samband mellan arbetsminne och lexikon påvisades hos barnen med CI samt hos kontrollgruppen. 
Inget samband kunde påvisas mellan undersökta bakgrundsvariabler och testresultat.
Denna uppsats undersöker hur den svenska modellen har influerat det svenska samhället under första halvan av 1900-talet och hur det var att leva under dess inflytande på 1960-talet. 
Under 60-talet dominerades det svenska samhället av de lagar och reformer som skapats av Socialdemokratiska Arbetarepartiet, SAP. 
Målet var att bygga upp Per Albin Hanssons vision av välfärdssamhället. 
Från det att han presenterade sin idé 1928, till och med 60-talet, genomgick Sverige en förvandling från ett agrart samhälle till ett industrialiserat. 
I vår analys av det svenska samhället under den här tidsperioden har vi använt oss av ett flertal konsumtionsteorier samt fokuserat på Raymond Williams tolkning av hegemonibegreppet. 
Hegemoni är ett organiskt begrepp som symboliserar den konsensus som råder inom ett samhälle vid en given tidpunkt. 
Efter att ha målat upp en bild av samhället och genomfört en förberedande analys har vi gått vidare med vår filmanalys för att studera hur det faktiska svenska samhället representeras i filmer från sin samtid. 
Vi har analyserat filmerna; Änglar, finns dom...? , Raggargänget och Sten Stensson kommer tillbaka. 
I analysen har vi lagt fokus på aspekter såsom kön, ålder och produktplacering. 
Vi har kommit fram till att filmerna i fråga presenterar en korrekt bild av det svenska samhället, det vill säga en så korrekt bild en film kan visa av ett samhälle utan att ha dokumentära intentioner. 
Vi har kommit till denna konklusion då miljöerna och normerna som existerade i det svenska samhället vid denna tidpunkt presenteras på ett korrekt sätt. 
Vi har också kommit till slutsatsen att även om produktplacering förekommer i filmerna, är detta främst i syftet att skapa en autentisk miljö.
Mariannes entusiastiska person som jag fick glädjen att möta och ta del av, löper som en gyllene tråd genom det här arbetet som jag vill delge er. 
Att Mariannes speciella och unika personlighet kommer fram på det sätt som det gör, beror mycket på valet av metod. 
Metoden bygger på att man får ta del av en person på ett djupare plan- en livsberättelse. 
Syftet att skriva om detta ämne är för det är viktigt hur jag som pedagog kan upptäcka de barn som far illa, eftersom barnen tillbringar den största delen av sin vakna tid i skolan. 
Arbetet handlar om hur jag som pedagog kan se/upptäcka barn som inte mår bra. 
Jag fick ett svar men det kom inte fram på det sättet jag räknade med. 
Svaret jag istället möttes av var inlindade i Mariannes engagerade berättelse om sitt liv som pedagog och människa. 
Jag möttes av en människa vars uppväxt var präglad av kärlek och omtanke som hon senare tagit med sig i sin pedagogik under 40 år. 
Att vara genuint intresserad av människor, men framför allt av barn har skapat den altruistiska pedagogen. 
Genom att ställa min litteratur bredvid Mariannes berättelse stod det klart för mig att sättet att upptäcka barn som far illa är att vara en besjälad pedagog.
Syftet med det här arbetet är att få en insyn i vad förskolebarn har för tankar om de frågor som berör döden.
Frågeställningen som besvaras är: "Vad har förskolebarn för tankar om döden?"
Kvalitativa intervjuer har skett med tio förskolebarn i åldrarna fyra till sex år vilka ligger till grund för undersökningen i arbetet. 
Även teckningar av barnen som förtydligar deras tankar ingår i undersökningen. 
Förskolebarnen tillhör samma förskola i Värmland.
Det som sägs i intervjuerna kan inte generaliseras att gälla alla förskolebarn, utan gäller enbart för de förskolebarn som intervjuerna är utförda med.
Undersökningsresultatet påvisar att förskolebarn har en öppen syn på döden. 
Barnen har haft tankar om det mesta som berör ämnet. 
Deras teckningar visade också en bred variation av tolkningar av döden.
Denna uppsats undersöker hur en utveckling av en medial identitet går till. 
Vilka faktorer får en medieidentitet att ändra dess mediala bild och framtoning? För att besvara denna fråga studerar jag en artistkarriär som har genomgått stora förändringar, vilka har inneburit att även dess medieidentitet kraftigt förändrat framtoning. 
Artistkarriären jag har valt att studera närmare är förgrundsfiguren från Latin Kings, Douglas "Dogge" Leóns. 
Metoden för att genomföra denna studie grundar sig i textanalys av de mediala framträdanden Dogge gjort i sin karriär.
Bakgrund:
Under 2000-talets början uppdagades ett antal företagsbedrägeriskandaler. 
Till följd av dem började investerare att ställa allt högre krav på företagens styrelser. 
I Sverige tog kodgruppen därför fram svensk kod för bolagsstyrning. 
Enligt koden för svenskbolagsstyrning är syftet "att förbättra styrningen av svenska bolag och ska utgöra god sed för bolagsstyrning". 
Tom Berggren som är medlem i svenska iskkapitalföreningen anser att ett av de största problemen som finns för att svenska IT-företag skall nå framgång, är bristen på kompetens och ambition.
Frågeställning:
Författaren har valt att definiera kompetens som utbildningsnivån för den enskilda styrelseledamoten. 
Yrkeserfarenhet som antalet år ledamoten har varit verksam i företagets styrelse. 
Engagemang definieras som antalet styrelser som den enskilda styrelseledamoten är verksam inom. 
Det skapade följande frågeställning:
Påverkar företagsstyrelsens kompetens, erfarenhet och engagemang svenska IT-företagets årliga resultat?
Syfte:
Uppsatsens syfte är att fastställa om det finns något samband mellan företagsstyrelsens sammansättning och nyckeltalet EVA i svenska IT-företag.
Metod:
En kvantitativ undersökning har genomförts med årsredovisningar som det huvudsakliga datamaterialet. 
Uppgifter om styrelseledamöterna samt underlag för beräkningarna av EVA-värden kommer ifrån respektive företags årsredovisning. 
En kvalitativ undersökning i form av en intervju har även ägt rum för diskussion av studiens resultat.
Slutsatser:
Styrelsen hos svenska IT-företag har en god kompetens, erfarenhet och är engagerade i sitt styrelsearbete. 
De är akademiskt utbildade och statistiskt sett har de en jämn fördelning mellan kandidat och magisterexamens. 
Det finns ett samband mellan styrelseledamöternas kompetens och företagets EVA-värde. 
Det finns däremot inget samband mellan nyckeltalet EVA och erfarenhet samt engagemang.
Orofaciala funktioner såsom mimik, tal, tuggning och sväljning är viktiga för livskvaliteten. 
Det råder generell brist på normerade test som bedömer dessa funktioner och därför har Nordiskt Orofacialt Test – Screening (NOT-S) utvecklats. 
Syftet med föreliggande studie var att normera NOT-S för barn med typisk utveckling i åldrarna 3:0-6:0 år. 
Testet består av en strukturerad intervjudel och en undersökningsdel med sex avsnitt vardera. 
Kalibrering utfördes innan testningen inleddes och visade på hög inter- och intrabedömaröverensstämmelse (94% respektive 96-99%). 
Det var 132 barn, 62 pojkar och 70 flickor, som deltog i testningen vilken utfördes på barnens förskolor. 
Resultatet visade att barn med typisk utveckling i åldersgruppen 3:0-3:11 år kan förväntas få en totalpoäng på 1,41 ± 0,96, barn i åldersgruppen 4:0-4:11 år en totalpoäng på 1,31 ± 1,04 samt barn i åldersgruppen 5:0-6:0 år en totalpoäng på 1,41 ± 0,94. 
Det fanns inga generella signifikanta ålders- eller könsskillnader. 
Signifikanta skillnader återfanns på enstaka frågor och uppgifter inom avsnitten Dregling (V), Näsandning (2) och Oral motorik (5). 
Sammanfattningsvis kan konstateras att NOT-S är ett lättadministrerat orofacialt test som med tillägg av denna normering har potential att bli ett välanvänt screeningmaterial för yrkesgrupper involverade vid bedömning av barns orofaciala funktion.
Syftet med examensarbetet har varit att undersöka möjligheterna att utveckla, producera och lansera en ny universell laddare. 
Målet har varit att kunna ladda så många modeller av så många produkter som möjligt, vilket innefattar mobiltelefoner, kameror, datorer och MP3-spelare etc. 
Arbetet skulle leda fram till ett förslag på produkt.
Genom att undersöka befintliga patent och produkter, har marknaden granskats och slutsatsen är att det finns en uppsjö av universella laddare på marknaden. 
Dock finns det få produkter som inger säkerhet, möjliggör multipel laddning och som är stationära. 
Dessa egenskaper blev grundstenar i den kravspecifikation som utarbetades. 
Genom en teknisk analys och kundundersökning sammanställdes ytterligare viktiga parametrar.
Resultatet blev en stationär produkt som kan ladda både en bärbar dator och flera mindre elektroniska produkter. 
Genom att använda en metod som i rapporten betecknas tappteknik kan rätt laddningsförhållande garanteras. 
Med hjälp av en mikroprocessor och produktspecifika tappar eller ändadaptrar kan laddning av i princip alla sorters produkter och modeller ske.
Arbetet har även innefattat konstruktion, CAD och prototypframtagning.
Vårt intresse för verksamhets- och systemutveckling har växt fram under vår studietid, då vi fått kunskap om att en av utvecklingstyperna har en mer prioriterad roll vid ett utvecklingsarbete. 
Efter att ha läst en del artiklar blev vi även intresserade av att jämföra vilka faktorer samt vem som är beslutstagare vid utveckling av organisationer i den statliga och privata sektorn. 
Detta för att se vilka eventuella skillnader respektive likheter det finns mellan dem.
Syftet med denna studie är att hitta de faktorer som är avgörande vid val att prioritera verksamhetsutveckling respektive systemutveckling. 
Samt att skapa en djupare förståelse för en organisations tänkande vid utveckling och hur utvecklingen skall genomföras.
Vi valde i denna studie att genomföra en kvalitativ studie där vi började med att tillägna oss relevant teori som förklarar och fördjupar läsaren i vad verksamhets- och systemutveckling är. 
Vidare utformade vi intervjufrågor utifrån vår problemformulering. 
Intervjufrågorna skickade vi ut till olika organisationer inom både den statliga och privata sektorn i Jönköpings län.
Utifrån den teori vi tillägnat oss och de svar vi fick in vid intervjuerna genomförde vi en analys som vi sedan kunde dra slutsatser från. 
Slutsatserna består av de faktorer som vi önskade få fram genom denna studie och presenteras i en matris.
Detta för att det ska vara lättare för läsaren att få en överblick över våra slutsatser. 
Genom matrisens uppbyggnad besvarar den vår problemformulering väldigt bra. 
Matrisen är uppbyggd enligt följande, den delar upp organisationerna i de två förut nämnda kategorierna, privat och statlig. 
Den skiljer även på faktorer för verksamhets- och systemutveckling samt vem som är beslutstagare.
Med beredning avses här den planering som görs för att möjliggöra och bestämma hur bearbetning skall utföras vid tillverkning av en enskild artikel. 
Med beredning avses även resultatet av ett beredningsarbete, vilket är en beskrivning av hur produktion skall utföras. 
Syftet med denna typ av beredning är att få vetskap om hur man tillverkar artikeln för effektivast produktion samt stödja konstruktörens arbete med att produktionsanpassa artikeln. 
Här återges mitt examensarbete med framtagning av förslag till en överskådlig grafisk framställning av beredningsarbetet på företaget Scania.
Scania har sedan tidigare en beskrivning för hur det inom företaget skall arbetas med beredning. 
Beskrivningen går under namnet 'Beredning för Bearbetning och Plåtformning, Arbetsmodell för Scania', men även kallad MPP (Machining Preparation Process). 
Scanias önskan är att komplettera arbetsmodellen med en Astrakanmodellerad grafisk beskrivning.
Astrakanmodellering är en metod och ett språk för att skapa verksamhetsmodeller. 
Astrakanmodelleringsspråket har tydligt släktskap med andra modelleringsspråk. 
Särskiljande för Astrakan är huvudidén att metoden ska vara ett hjälpmedel för att på ett enkelt sätt beskriva en verksamhet. 
Metodens förvaltare har dokumenterat metoden kortfattat. 
Dess notation och regelverk är mindre utförliga relativt närbesläktade språk.
Den grafiska beskrivningen presenteras som en processmodell för beredning. 
För att uppnå målet att den grafiska beskrivningen skall vara överskådlig och samtidigt vara så entydig som möjligt så kompletteras den med två begreppsmodeller. 
Det är en modell för beredningstekniska begrepp och en modell för modelleringsspråkliga begrepp. 
Modellerna definierar viktiga begrepp och skall användas som stöd för att tolka processmodellen för beredning som avsett.
Syftet med Processmodellen för beredning är att beskriva hur beredning skall utföras. 
Synvinkel för modellen är en beredare eller annan person som arbetar med beredning. 
Processmodellen är uppdelad i delprocesser och kan presenteras och läsas i olika detaljeringsgrad. 
Processmodellen har beredningen som förädlingsobjekt. 
Den beredning som beskriver hur produktionen skall utföras.
Examensarbetet har konkret resulterat i tre modeller som kan användas som komplement till tidigare beskrivning av beredningsarbete på Scania. 
Modellerna ger ett processorienterat modellperspektiv på arbetsmodellen för beredning på Scania. 
Arbetet har även gett mig och arbetsgruppen för MPP arbetsmodell en ökad kunskap och förståelse kring modellering och tolkning av modeller.
Under många år har opinionsbildare såsom Mäklarsamfundet arbetat för en förnyelse av Fastighetsmäklarlagen.
Den 31 december 2007 skall utredningsarbetet kring den nya Fastighetsmäklarlagen vara klart och en av de frågor som utredningsgruppen avhandlar är huruvida fastighetsmäklare skall få förmedla kringtjänster till sina kunder eller ej. 
Mot bakgrund till det utredningsarbete som för närvarande förs kring den nya Fastighetsmäklarlagen har det varit mitt syfte med denna promemoria att beskriva komplexiteten om kringtjänsternas vara eller icke vara, och med vilken nytta tjänsten kan bidra med till konsumenterna och fastighetsmäklarbranschen. 
Jag har under mitt arbete stött på teorimotsättningar då den ena teorin förespråkar att det är kunden som är i fokus och bestämmer, menar den andra teorin att det är ej bra att ha en alltför spridd tjänst då tjänsteföretaget skall fokusera på kärntjänsten. 
När dessa teorier har sammanvävts med empirin anser jag att fastighetsmäklarföretagen kan använda sig av kringtjänsterna för att positionera sig gentemot sina konkurrenter och framförallt för mindre fastighetsbyråer kan det vara avgörande för hur de skall överleva i framtiden.
Sammanfattning
Vår värld står inför nya utmaningar i form av ett förändrat klimat. 
FN: s klimatpanel har fastslagit att det är människan som bär det största ansvaret, men också att vi kan begränsa verkningarna genom att förändra vår livsstil. 
Detta kräver att information når ut till människor vilket i praktiken innebär att skolan måste arbeta med dessa frågor. 
Det betyder också att lärarna måste vara medvetna och ge frågorna det utrymme som behövs. 
Syftet är att se om denna medvetenhet finns idag, bland aktiva lärare och lärarstudenter, och om synsättet skiljer sig åt mellan dem, men också om deras uppfattningar är i paritet till kursplanen. 
För att ta reda på det har jag formulerat tre forskningsfrågor: 
Vilken uppfattning av geografiämnet har lärarstudenter, inom geografiämnet vid karlstads universitet, och vilken vikt lägger de vid miljöfrågor? 
Vilken uppfattning av geografiämnet har behöriga aktiva lärare och vilken vikt lägger de vid miljöfrågor? 
Föreligger det någon skillnad mellan aktiva lärare och lärarstudenter gällande uppfattningar om geografiämnet? 
I syfte till att besvara forskningsfrågorna har jag använt mig av en kvalitativ metod i form av intervjuer vilka analyseras utifrån en tematisk innehållsanalys. 
Resultatet visar att båda urvalsgrupperna lägger stor vikt vid miljöfrågor i undervisningen med viss övervikt för lärarstudenterna. 
I övrigt uppfattar urvalsgrupperna geografiämnet i paritet med de rådande kursplanerna, förutom något undantag för respektive intervjuobjekt. 
Slutsatsen blir att miljöfrågor uppfattas som en viktig del i geografiämnet, lärarstudenterna uppfattar kulturgeografin som en viktigare del i geografiämnet än vad de aktiva lärarna gör medan det är tvärtom gällande kart/namn/platsgeografi. 
Vidare framkommer att endogena (inre)och exogena (yttre) krafter får den största svarsfrekvensen gällande uppfattningarna av geografiämnet.
Idag bedrivs en stor del av forskningen vid högskolor och universitet i projektform. 
Detta gäller inte minst inom teknik, naturvetenskap och medicin, men numer också inom samhällsvetenskap.
Det är vanligt att olika personalkategorier så som exempelvis professorer,docenter, och doktorander ingår i projekten. 
Projektledaren är oftast den som har ansökt om projektmedlen, eller den person som är mest vetenskapligt meriterad vid avdelningen, vilket ofta är en professor eller docent med lång erfarenhet. 
Av de här personerna förväntar sig organisationen ofta underverk. 
De ska medverka i alla möjliga typer av aktiviteter, som exempelvis handledning av doktorander,undervisning, medverkande vid och organiserande av konferenser,ansökan om medel för nya projekt och vara avdelningens ansikte utåt. 
Dessutom ska de också agera projektledare för en eller flera parallella projekt.
I den här uppsatsen redovisar vi först en kartläggning av projektledarkompetens hos projektledare i forskningsprojekt vid Karlstads universitet. 
Kartläggningen har gjorts med stöd av två enkätundersökningar och sex stycken kompletterande intervjuer. 
Såväl professorer och docenter som doktorander har medverkat i studien. 
Kartläggningen visar klart och tydligt att de flesta projektledarna leder projekten baserat på tidigare erfarenheter och merparten saknar ledarskapsutbildning. 
Detta innebär att beprövade projektledningsmetoder och tekniker sällan används.
Baserat på resultat från enkätundersökningarna, intervjuerna och deltagande observationer presenterar vi dessutom fyra konkreta förbättringsåtgärder för forskningsprojekt vid Karlstads universitet. 
Åtgärderna tror vi kan effektivisera forskningsprojekten och därmed medföra en besparing för Karlstads universitet. 
Den första åtgärden är att utveckla en kurs i projektledningsmetodik, som sedan erbjuds till alla projektledare vid Karlstads universitet.
Den andra åtgärden är att bygga upp en eller flera erfarenhetsnätverk bland aktiva projektledare. 
Den tredje åtgärden är att skapa ett mentorsprogram för stöd åt nya projektledare. 
Den fjärde och sista åtgärden är att etablera en grupp med erfarna projektledare som kan ge stöd åt andra projektledare.
Internkommunikation är av mycket stor vikt för en organisations framgång. 
Landstinget i Värmland är en stor organisation med många mellanchefer på olika befattningar. 
Alla dessa får varje vecka ett mail om att ett nytt chefsbrev, Chef, utkommit på intranätet. 
Med min uppsats undersöker jag hur cheferna uppfattar och använder sig av detta chefsbrev samt om uppfattning och användning skiljer sig åt bland olika befattningsgrupper. 
Jag önskar ta reda på om Chef behövs som en del av landstingets interna kommunikation.
Studiens frågeställningar försöker jag besvara genom att använda mig av en kvantitativ metod i form av en enkät som skickas ut till alla mottagare av chefsbrevet. 
Resultatet av studien visar att Chef till stor del verkar vara en lyckad informationskanal. 
En majoritet av cheferna tittar igenom åtminstone de flesta numren, anser att en större del av innehållet känns viktigt att ta del av och anser inte att någon annan kanal skulle kunna ersätta chefsbrevet. 
Majoriteten upplever också att innehållet är aktuellt och tillförlitligt samt att de har ganska stor nytta av brevet i sitt arbete.
Ett uttalat syfte med Chef är att cheferna i Landstinget i Värmland ska läsa det och vidareinformera till sina medarbetare. 
Resultatet visar att en majoritet av cheferna ofta vidareinformerar men jag anser att den andel som inte gör det är alltför stor. 
Chefernas kommunikativa ansvar bör därför tydligare beskrivas så att de förstår vad som förväntas av dem, samtidigt som de bör få hjälp att utveckla sin kommunikativa förmåga.
Skillnaderna mellan hur de olika befattningsgrupperna uppfattar och använder sig av Chef är inte så stora men vissa skillnader finns. 
Divisionscheferna som befinner sig högt upp på organisationsschemat och ingår i en ledningsgrupp är mer nöjda med Chef än vad avdelningschefer och chefer inom serviceverksamheter, som befinner sig längre ifrån ledningen är. 
Ansvariga bör fundera på hur dessa skillnader skulle kunna minskas.
De problem som visat sig finnas bör åtgärdas men är givetvis inte anledning nog att avveckla chefsbrevet, som ändå är en väl fungerande, etablerad kanal. 
Det visar sig alltså att en bra Chef går hem.
Pliktverket genomförde under 2006 en stor förändring för att spara 100 miljoner kronor.
Resultatet blev att 131 medarbetare sades upp och två regionkontor lades ner. 
Syftet med denna uppsats är att undersöka anledningarna till negativa omdömen om Pliktverkets interna kommunikation under förändringsprocessen 2006 och komma fram till lösningsförslag på de bakomliggande problemen så att den interna kommunikationen kan utvecklas.
Kommunikation under förändring är ett stort område och därför har jag valt att begränsa mig till fyra områden som Pliktverket i en enkätundersökning funnit att det varit problem med.
Jag har arbetat utifrån följande problemområden:
Tillförlitlighet – Har tillförlitligheten till processen och informationen påverkats av problemen med kommunikationen?
Förväntningar – Har Pliktverket skapat orimliga förväntningar på förändringsarbetet via medarbetarutbildning?
Delaktighet – Varför får delaktigheten lågt betyg och hur har medarbetarna varit delaktiga?
Dialog – Varför får dialogen under processen dåligt betyg?
Samtalsintervjuer med medarbetare vid Pliktverkets kvarvarande regionkontor och huvudkontoret har använts som metod.
Jag har bland annat kunnat dra följande slutsatser:
- Förändringen har varit toppstyrd utan delaktighet för medarbetarna
- Monolog har förekommit istället för dialog, vilket har lett till att tillförlitligheten och förtroendet för processen har blivit lågt.
- Delaktigheten inom organisationen har av allt att döma varit dålig redan innan förändringsprocessen.
- Medarbetarutbildningen som genomförts tidigare har gett medarbetarna förväntningar på att få vara delaktiga under en förändringsprocess.
- Dålig tillgänglighet till ansvariga och chefer har gjort att dialogen blivit dålig.
- Förändringens syfte är dåligt förankrad i organisationen på grund av dålig dialog.
En allt mer föränderlig marknad har medfört en ökad konkurrens och förändrade förutsättningar för dagens företag. 
De ökade kraven från marknaden har gjort att synen på företagens styrning har förändrats och en mer processinriktad och kundanpassad verksamhetsstyrning har de senaste åren presenterats i litteratur och studier. 
Företagens ekonomistyrning i praktiken har däremot inte utvecklats i samma takt som dessa nya idéer. 
Denna kvalitativa studies syfte är att undersöka och analysera de faktorer som kan hindra eller försvåra en utveckling av ett företags ekonomistyrning. 
Controllers och ekonomichefer har intervjuats för att undersöka på vilket sätt deras ekonomifunktioners rutiner, struktur och resurser påverkar möjligheten att utveckla företagets ekonomistyrning mot en mer horisontellt riktad verksamhetsstyrning. 
Studien visar att ekonomisystemen är uppbyggda av fasta rutiner och regler. 
Detta medför att de tar lång tid att förändra eftersom de blivit rotade i företagets organisationsstruktur och utgör en trygghet för företagets anställda. 
Undersökningen visar även att ekonomifunktionens resurser inte i sig är något hinder mot en fortsatt utveckling av företagets styrning, så länge det går att motivera att en investering ger resultat visar studien att det ofta finnas möjlighet till nya satsningar. 
Snarare tyder det mesta på att det är controllerns förmåga och vilja att identifiera att det behövs en förändring som är det största hindret mot en utveckling av företagets ekonomistyrning.
Avsikten med studien är att undersöka relationen mellan valberedning, ägare och styrelse samt utifrån detta studera vilken roll valberedningen har, enligt den Svenska Koden.
Vi har utgått ifrån en deduktiv ansats, där vi både har genomfört en kvantitativ och en kvalitativ undersökning. 
Den kvalitativa studien baseras på djupintervjuer av ledamöter i svenska börsnoterade företag, medan den kvantitativa undersökningen resulterar i en statistisk undersökning, som utgår från bolagsstyrningsrapporter i årsredovisningar från 2006.
I det teoretiska perspektivet tas den Svenska Koden för bolagsstyrning upp som utgångspunkt och kompletteras med Aktiebolagsslagen (ABL), agentteorin, intressentmodellen, coporate governance, CSR-modellen samt ett genusperspektiv.
I empirin redovisas respondenternas yttranden samt den statistiska undersökningen.
Vi har med hjälp av empiri och analys kommit fram till ett antal slutsatser; valberedningen har endast en uppgift, vilken är att ta fram förslag om nya ledamöter till styrelsen. 
Förslagen ska leda till att styrelsen får en så bra sammansättning som möjligt. 
Valberedningen har till viss del ökat förtroendet för bolagen, genom att processen blivit tydligare samt mer transparant. 
Vår undersökning visar att nästan samtliga företag som är noterade på Stockholmsbörsens LargeCap-lista, använder sig av en valberedning, vilket vi ser som ett bra tecken. 
Koden är fortfarande relativt ny och är därför ännu inte fulländad. 
Koden är även unik i ett internationellt perspektiv och den svenska företagskulturen verkar anpassa sig efter Kodens riktlinjer.
Grunden med kalkylering är att skapa en logisk modell som avspeglar ett företags relevanta kostnadsmekanismer. 
På 1980-talet växte ABC-kalkylen fram pga. företagens nya sätt att arbeta på t.ex. genom användning av ny teknik, kundanpassning, kvalitetssatsning och produktdifferentiering. 
Hur omkostnaderna ska kalkyleras rättvist enligt ABC-metoden har varit en omdebatterad fråga ända sedan kalkylmetoden uppstod.
Idén med uppsatsen uppkom i januari 2007 under en diskussion med det svenska stålföretaget Uddeholm Tooling AB där vi kom fram till att det vore intressant att undersöka fördelningen av företagets omkostnader.
Syftet med uppsatsen är att undersöka om omkostnaderna kan fördelas på respektive produkt och se om Uddeholm Tooling AB:s tumregel är den mest lämpliga metoden för företaget. 
Uddeholm Tooling AB fördelar inte försäljnings-, lager- och administrationsomkostnader direkt ner i självkostnaden.
Metodvalet för undersökningen är en kvalitativ fallstudie med en deduktiv ansats. 
För att genomföra undersökningen valde vi tillsammans med Uddeholm Tooling AB ut tre produkter som representerar tre olika tillverkningskostnader samt att vi intervjuade representanter för försäljnings-, logistik-, lager- och ekonomiavdelningen.
Med hjälp av vårt framarbetade material kan vi i vår slutsats konstatera att den nuvarande kalkyleringsmetoden som Uddeholm Tooling AB använder sig av är den mest lämpade arbetsmetoden för företaget. 
I nuläget är det svårt att avgöra om omkostnaderna kan fördelas rättvist på produkterna, eftersom de anställda på respektive avdelning för de undersökta omkostnaderna inte har en arbetsfördelning på produkterna. 
Dock har vi lyckats att konstatera att det skiljer i arbetsbörda i själva lagerhanteringen, som därav skulle kunna härledas till respektive produkt. 
Resultatet av vår studie visar dock att företagets arbetssätt inte utförs enligt en logisk modell som avspeglar företagets relevanta kostnadsmekanismer pga. företagets tumregel. 
Arbetssättet visar ändå att kalkyleringsmetoden är praktiskt användbar i det dagliga arbetet.
Utvecklingen inom redovisningsområdet har gått i mycket rask takt. 
Den svenska lagstiftningen har anpassats till EG-rätten och gjort redovisningen onödigt svår och komplicerad för onoterade svenska företag. 
På grund av detta har bokföringsnämnden idag delat upp företag i fyra olika kategorier med olika redovisningskrav beroende på storlek. 
Dessa kategorier benämns K1, K2, K3 och K4. 
Denna kandidatuppsats är begränsad till att enbart behandla K3.
Bokföringsnämnden har än så länge enbart lagt fram ett utkast för K3-regelverket.
Informationen i utkastet är så pass tunn att syftet med uppsatsen är att försöka ta reda på hur det nya regelverket bör utformas, så att det gynnar så många företag som möjligt inom denna kategori. 
I teorin beskrivs till en början de regler som gäller för företag idag, i väntan på att det nya regelverket.
Teorin avslutas med en övergripande beskrivning av K3-regelverket men även en härledning från utkastet till Redovisningsrådets rekommendationer.
Empirin har framställts genom kvalitativ metod där vi via intervjuer med revisorer i Karlstad diskuterat kring hur det nya K3-regelverket bör se ut och kan tänkas påverka de företag som hamnar inom K3.
Efter att ha analyserat empirin och teorin kan det konstateras att många företag hamnar inom K3. 
En del är tidigare medelstora företag enligt de gamla gränsvärdena och dessa företag kommer troligtvis att få försvårade regler. 
De större K3-företagen kan däremot få förenklade regler då det nya regelverket kommer att innehålla mindre tilläggsupplysningar än dagens regler. 
Vi anser att det är svårt att lösa denna problematik utan att riva den struktur som finns inom K3. 
Vår slutsats är att de mindre K3-företagen bör ha mindre krav med undantagsregler än om man jämför med de större K3-företagen då det i de mindre K3-företagen inte finns ett speciellt stort externt intresse.
Älgen är en viktig art, både ekonomiskt och ekologiskt, och all kunskap är viktig för att även i framtiden kunna sköta en sund älgstam. 
Trots flertalet studier finns det många frågetecken om älgens habitatval i Sverige. 
En ökad exploateringstakt och nya infrastrukturprojekt hotar att fragmentera och isolera populationer av älg. 
Habitatvalet hos 22 älgar, 8 tjurar och 14 kor, i sydvästra Sverige studerades mellan februari 2002 och december 2005. 
Älgarna sövdes och utrustades med GPS-sändare, deras positioner registrerades varannan timma och det totala antalet positioner under den 46 månader långa studietiden var 71103 stycken. 
Data från varje älg delades in i 4 säsonger; vår, sommar, höst och vinter, baserat på klimat och älgens biologi. 
Totalt genererades 125 hemområden baserade på säsong, och valet av habitat inom varje hemområde studerades med hjälp av Euclidean distance-based analysis. 
En omklassificerad digital marktäckedata användes som var indelad i 6 olika klasser; odlad mark, hygge, barrskog, lövskog, myrmark och berg i dagen. 
Resultaten visade att det var skillnad mellan könen i hur de väljer habitat. 
Tjurarna var signifikant närmare barrskog och hyggen än korna, men både tjurar och kor selekterade för hyggen och undvek odlad mark inom deras hemområden.
Undersökningens syfte är att studera hur anställda i kunskapsföretag utvecklar kompetens för att klara det dagliga arbetet Fokus ligger på den informella kompetensutvecklingen. 
De teoretiska utgångspunkterna innefattar teorier om lärande och kompetensutveckling, organisationsförändring och utvärdering samt professionell reflektion. 
I undersökningen används narrativ analys och intervjuer vilket baseras på uppfattningen att kunskap om verkligheten bara kan nås genom språk och kommunikation.
De postmoderna uppfattningarna om den snabba (tekniska) utvecklingen och kravet på att vara uppdaterad påverkar starkt informanternas syn på arbetslivet, liksom känslan av att inte ha tillräckligt med tid för all den kompetensutveckling som önskas. 
Men tiden arbetar också för kompetensen eftersom erfarenhet är något som utvecklas över tid. 
Resultaten leder fram till slutsatsen att både drivkrafterna till och målet för kompetensutveckling är att skapa en begriplig och hanterbar verklighet.
Våra kyrkor är en viktig del av samhället, och är en kulturskatt som måste vårdas. 
Kyrkorna använder dock väldigt mycket energi till uppvärmning varje år. 
Detta beror på att de flesta av dem är gamla och att energieffektivitet ej varit en prioriterad fråga i deras verksamhet. 
Grinstad kyrka är en kyrka med hög energianvändning som trots att den endast är uppvärmd vid förrättningar använder lika mycket energi som två medelvillor. 
Kyrkan är från 1200-talet, är byggd i tegel och värms idag upp av en oljepanna i ett vattenburet system samt några elradiatorer. 
Det finns planer på att byta ut oljepannan mot närvärme.
Syftet med examensarbetet var att undersöka och ge församlingen en inblick i vart den energi som tillförs kyrkan tar vägen, hur mängden tillförd energi kan minskas genom energieffektiviseringsåtgärder samt vilken miljöpåverkan värmekällan i dagens uppvärmningssystem har jämfört med värmekällan i det planerade närvärmenätet.
Målet var att svara på följande frågor:
- Var sker de största energiförlusterna i kyrkan och hur skall dessa kunna minskas genom energieffektiviseringsåtgärder?
- Hur skall kyrkans värmesystem dimensioneras med avseende på kyrkans värmeeffektbehov?
- Hur skulle miljöpåverkan till följd av kyrkans uppvärmning förändras vid anslutning till det planerade närvärmenätet.
Det värmesystem som ansågs passa Grinstad kyrka bäst var ett vattenburet värmesystem som värmer kyrkan intermittent. 
Det ansågs även lämpligt att värma upp på 6 timmar från en grundtemperatur av 8°C till en förrättningstemperatur av 18°C. 
Värmesystemet måste då ha effekten 22,5 kW, vilket är en effekt som är högre än dagens system kan avge. 
Därför gavs förslaget att komplettera dagens system med kamflänsrör under några av kyrkbänkarna.
De största energiförlusterna i kyrkan visade sig vara genom taket och genom att isolera detta kan förlusterna genom det minskas med 85 %. 
Grundtemperaturen i kyrkan är idag högre än vad som behövs och genom att sänka den 4ºC kan energianvändningen för grundvärmen minskas med 18 %.
Bytet från en central oljepanna till biobränsleeldad närvärme skulle leda till att utsläppen av koldioxid och svavel att minska, medan utsläppen från stoft, koloxid och svavel kommer att öka.
Denna rapport omfattar ett 15 poängs (22,5 högskolepoäng) examensarbete vid Karlstads universitet. 
Arbetet har utförts på plats hos BAE Systems Bofors i Karlskoga. 
Företaget ville kunna styra en radiostyrd leksaksstridsvagn med en laserpekare. 
En kamera ansluten till en digital signalprocessor (DSP) skulle kunna detektera var en laserpunkt befinner sig och styra stridsvagnen mot den.
Ett styrgränssnitt mellan DSP:n och leksaksstridsvagnen konstruerades och byggdes med hjälp av en programmerbar logisk krets. 
Leksaksstridsvagnens interna signalsystem analyserades. 
En manchesterkodad signal i form av ett 32-bitars seriellt kodord hittades, vilket ursprungligen kom från radiostyrningen. 
Ett styrgränssnitt konstruerades kring en CPLD (Complex Programmable Logic Device) vilken programmerades med VHDL (Very high speed integrated Hardware Description Language) som återskapar den Manchesterkodade styrsignalen.
Gränssnittet ansluter till DSP:n som kontrollerar stridsvagnens styrning och övriga funktioner till fullo. 
Kommunikationen mellan styrgränssnittet och DSP:n sker via ett parallellgränssnitt som är 16-bitar brett. 
13 bitar är datasignaler och övriga tre är "styrbitar" som konfigurerar gränssnittet. 
En applikation integrerades i projektet för att demonstrera styrgränssnittets funktion. 
DSP:n tolkar var en laserpunkt befinner sig inom ett kameraområde och skickar motsvarande styrsignaler till leksaksstridsvagnen.
Syftet med denna undersökning har varit att beskriva och analysera sex pedagogers syn på sitt ledarskap. 
För att göra detta har jag genomfört sex kvalitativa intervjuer med olika pedagoger. 
De intervjuade är: tre förskolelärare, två lärare för yngre barn och en fritidspedagog. 
Pedagogerna är från olika städer och olika arbetslag. 
Jag har utfört undersökningen utifrån fyra huvudfrågor:
- Vad innebär ledarskapet?
- Vad är det som påverkar ledarskapet?
- Hur kan man utveckla sig själv som ledare?
- Vilken sorts ledare behöver barn idag?
Resultatet visar att ledarskapet i läraryrket framförallt innebär att lära barnen det sociala samspelet. 
Pedagogerna anser att ledarskapet påverkas av en rad faktorer, bl.a. av barngruppen, kollegorna, den egna personligheten och egna erfarenheter. 
Utvecklingen till att bli en bättre ledare sker genom att man får erfarenhet. 
Man utvecklar sig själv bl.a. genom att pröva olika metoder och genom att lära av andra ledare. 
Intervjupersonerna anser att barn idag bl.a. behöver en tydlig ledare som kan sätta gränser och samtidigt vara en lyhörd ledare som lyssnar på barnen.
Syfte och frågeställningar
Syftet med studien är att undersöka förekomst, hantering och upplevda orsaker till mentala blockeringar inom kvinnlig truppgymnastik på nationell ungdoms- och juniornivå.
- Vilken typ av övning är den vanligaste mentala blockeringen inom kvinnlig truppgymnastik?
- Hur visar sig blockeringarna enligt gymnasterna och tränarna?
- Vilka orsaker till uppkomsten av mentala blockeringar kan utläsas utifrån gymnasterna och tränarnas berättelser?
- På vilka sätt har gymnaster och tränare försökt hantera mentala blockeringar?
Metod
Studien inleddes med en litteratursökning för att finna tidigare forskning. 
Därefter utformades en enkät i två versioner (för tränare och gymnaster) och dessa delades ut till gymnaster och tränare på nationell ungdoms- och juniornivå i sex olika föreningar. 
Gymnasterna valdes efter tränings- och tävlingsnivå och har en medelålder på 14 år.
Resultat
Resultatet visade att mentala blockeringar är ett mycket vanligt fenomen inom truppgymnastiken och något som majoriteten av gymnasterna någon gång drabbats av. 
Blockeringarna visar sig ofta genom att gymnasten vägrar eller helt utesluter övningen ur sin träning och blockeringarna är vanligast i grenen tumbling. 
Dock visade studien att de flesta gymnaster upplever blockeringar i mer än ett redskap. 
Volter som roterar baklänges tenderade att vara den typ av övning som flest gymnaster har blockeringar för.
Detta ansågs främst bero på att gymnasterna i fråga inte tror att de kommer att lyckas med övningen följt av orsaker som tidigare skador och mental omognad. 
De allra flesta gymnaster och tränare har på något sätt försökt behandla problemet, främst genom fysiska åtgärder och har i situationer med mentala blockeringar känt sig rädda, frustrerade och misslyckade.
Slutsats
Problematiken kring mentala blockeringar är stor och få gymnaster och tränare vet hur de kan hantera dessa.
Behovet av fortsatt forskning inom området samt större fokus på mental träning inom förbundets utbildningar är stort.
Den här rapporten handlar om det examensarbete som utförts mot Volvo 3P genom forskningsprojektet Viktor. 
Viktor är ett projekt som ska visa möjligheten med virtuell produktframtagning av gjutna komponenter. 
Volvo 3P är ett företag som utvecklar lastbilar. 
Uppgiften har varit att visa möjligheten att använda topologioptimering som ett verktyg i konstruktionsfasen. 
Detta har gjorts med hjälp av ett case som erhållits från Volvo 3P. 
Ett nytt koncept för en av deras lastbilsnav har tagits fram. 
Konceptet visar på högre styvhet och en lägre spänningsnivå än dagens originalnav. 
Konceptet hade förmodligen aldrig uppkommit om det inte hade varit för topologioptimeringen. 
Rapporten behandlar de steg som utförs vid en topologioptimering med programvaran Altair Hypermesh Optistruct. 
För att verifiera de resultat som erhållits från topologioptimeringen har koncepten analyserats i Abaqus. 
Rapporten tar även upp begränsningar och svårigheter som användaren kan komma att stöta på under arbetets gång.
Detta examensarbete handlar om drama som pedagogik, vad det är, hur man gör och varför man gör det. 
Mitt syfte med den här uppsatsen är att lyfta fram kunskap om hur vi pedagoger ska kunna hjälpa elever i våra klasser genom att använda drama som metod för kunskap och utveckling. 
Arbetet innefattar tre intervjuer samt litteraturstudier om ämnet. 
Individerna som jag har intervjuat är en klasslärare på mellanstadiet, en dramalärare samt en barnteaterförfattarinna. 
Intervjuerna innehöll frågor som rörde drama som pedagogik och hur de som pedagoger kommer i kontakt med detta, vad de tycker om drama som pedagogik, samt vad man kan använda det till och vilka fördelar som blir följden av användandet.
Jag kom fram till att drama som pedagogik är en metod med vilken elever och lärare lär sig mer om sig själva, varandra och världen. 
Jag kom också fram till att drama som pedagogik verkar både personlighetsutvecklande och grupputvecklande samtidigt som den hjälper eleverna på ett stimulerande, kreativt och roligt sätt mot sina kunskapsmål och är därför en bra metod. 
Jag kom också fram till att vi pedagoger genom att bjuda på oss själva, samtidigt som vi involverar eleverna i en beslutandeprocess om sitt eget lärande inom dramats ramar, där vi verkar som medagerare för att inspirera, stimulera och styra våra elever, så att de upplever att kunskapsinhämtande är roligt och intressant, utövar en givande pedagogik som stärker individerna i gruppen.
I min uppsats har jag valt att undersöka hur och i vilket syfte pedagoger använder sig av musik i förskol
an. 
Undersökningen baserar sig på litteratur och kvalitativa intervjuer. 
Fyra förskolelärare har intervjuats och resultatet visar att samtliga förskolelärare använder sig av musik med syfte att stimulera barnens språkliga, motoriska och sociala utveckling. 
Trots detta tycks musiken inte användas tillräckligt i förskolan. 
Det finns få situationer, där barnen själva spontant får skapa och experimentera med musik. 
Arbete med instrumenten fungerar dåligt,de finns inte tillgängliga för barnen mer än vid styrda aktiviteter som dessutom förekommer sällan. 
Undersökningen innehåller även en analys över orsakerna till detta.
Syfte
Syftet med föreliggande studie är att jämföra tre manliga elittränares arbetssätt i rollen som coach, analysera deras synsätt på coachrollen samt beskriva vägen till framgång.
Frågeställningar
Hur kan de tre elittränarnas bakgrund beskrivas?
På vilket sätt ser de tre elittränarna på sin roll som coach och hur arbetar de i praktiken?
Hur ser kollegorna och spelarna, i det egna laget, på elittränaren i rollen som coach?
Om det finns några gemensamma nämnare för tränarna, vilka är de?
Vilka är framgångsfaktorerna?
Metod
Undersökningen är genomförd i tre steg:
1. Observationer av de tre elittränarna i rollen som coach under en tävlingsmatch. 
Dessa obser-vationer är gjorda utifrån ett eget författat observationsprotokoll.
2. Halvstrukturerade intervjuer med en assisterande tränare och en lagkapten, inom respektive idrott, för att få deras syn på tränaren ifråga.
3. Halvstrukturerade intervjuer med de tre elittränarna.
Resultat
De undersökta tränarna har en tydlig självbild. 
Denna självbild förstärktes genom observatio-ner och kompletterande intervjuer. 
Alla intervjuade tilltalades av de aktuella tränarnas lugna coachstil. 
Tränarna är präglade av sin idrottsliga uppväxt, de har många av sina värderingar därifrån. 
De är kunniga och noggranna i sitt arbete och strävar efter att skapa en positiv och stimulerande miljö. 
Kommunikation är ett arbetsredskap.
Coacherna har många gemensamma nämnare, exempelvis: uppväxtmiljö, långa karriärer inom respektive idrott, engagemang, öd-mjukhet och situationsanpassat ledarskap.
Slutsats
De tre undersökta tränarna har i mångt och mycket samma arbetssätt. 
De sätter laget och den enskilde spelaren i fokus under såväl träning som match. 
Vid dessa tillfällen har tränarna total koncentration på laget och spelarna. 
De arbetar mycket hårt för att laget ska nå framgång. 
Vä-gen till framgång kan bero på tillfälligheter, men hårt arbete och ödmjukhet inför uppgiften, här och nu, ger troligtvis utslag i det långa loppet.
Nuvarande implementationer av distribuerade hashtabeller (DHT) har en begränsad storlek för data som kan lagras, som t.ex. OpenDHTs datastorleks gräns på 1kByte. 
Är det möjligt att lagra filer större än 1kByte med DHT-tekniken? Finns det någon lösning för att skydda de data som lagrats utan att försämra prestandan? Vår lösning var att utveckla en klient- och servermjukvara. 
Mjukvaran använder sig av DHT tekniken för att dela upp filer och distribuera delarna över ett serverkluster. 
För att se om mjukvaran fungerade som tänkt, gjorde vi ett test utifrån de inledande frågorna. 
Testet visade att det är möjligt att lagra filer större än 1kByte, säkert med DHT tekniken utan att förlora för mycket prestanda.
De allra flesta fastighetsmäklare i Sverige arbetar med provisionslön. 
Syftet med det här arbetet är därför att förhoppningsvis skapa en diskussion i fastighetsmäklarbranschen om det är nödvändigt med provisionslön. 
Vi har intervjuat sex fastighetsmäklare och bland annat kommit fram till att det är dags för en förändring i fastighetsmäklarbranschen och att det bör föras en gemensam diskussion om lönesättningen.
Sammandrag
Detta examensarbete bygger på en fallstudie av en manlig pedagog i förskolan. 
En aktuell fråga i dagens debatt är bristen på män i förskolan, vilket medför att en närmare granskning av manliga pedagoger kontra kvinnliga pedagoger är befogad. 
Frågan är på vilket sätt manliga pedagogers tänkande och beteende skiljer sig från kvinnliga pedagogers motsvarande? Syftet med den här undersökningen är att med hjälp av videoinspelning i detalj analysera en manlig pedagogs arbete tillsammans med barnen på en förskola. 
Speciellt söker jag vilka uppgifter en manlig pedagog väljer att utföra tillsammans med barnen, hur han väljer att utföra dem och vilket språk han använder. 
Den empiriska basen är observationer (videofilm) av en manlig pedagogs arbete under två dagar. 
Observationerna kompletterades även med en intervju för att genom den få en bredare bild och ett sammanhang utifrån respondentens perspektiv.
Undersökningen visar i sammanfattning att den manlige pedagogen skiljer sig i ganska hög grad från sina kvinnliga pedagoger och deras arbetssätt. 
När han valde aktiviteter själv prioriterade han att busa med barnen och själv leka barn. 
Han deltog i leken som en jämlik, medan den kvinnliga pedagogen behöll sin pedagogroll även i leken. 
Språkmässigt använder han sig av färre ord och även av en mer direkt kommunikation. 
Han ser sig själv som ett komplement i den kvinnodominerade pedagoggruppen. 
Genom att vara ett komplement ser han till att bidra med, enligt honom, typiskt manliga saker och aktiviteter.
Nyckelord: manlig pedagog, könsroller, manligt språk, förskolan.
C-uppsats vars huvudsyfte var att undersöka hur stor igenkänning människor har av företagsmärken utan att logotypen finns med. 
Genom att arbeta med både en kvalitativ och kvantitativ metod har vi fått fram våra resultat, detta genom att våra respondenter besvarade en enkät. 
Våra teoretiska perspektiv kommer från en blandning av olika ämnesområden, så som psykologi och informationsdesign med fördjupningar i bland annat perception, objektsigenkänning, symbolik och färgers betydelse. 
Genom våra undersökningar kom vi fram till att det inte finns något enkelt svar på huruvida märken känns igen eller inte. 
Bland våra utvalda märken var könsbundenheten låg, och ålder har viss betydelse för igenkänningen. 
Detta genom att äldre respondenter hade en högre igenkänning än de yngre.
Syftet med detta examensarbete var att undersöka möjligheten att använda en Dynamic Mechanic Thermal Analyzer (DMTA) för att mäta ökningen av styvhet som följd av filmbildning av latex i en torr bestrykning.
Två olika latexer användes för experimenten, en med Tg = 36°C (hård) och en med Tg = 8°C (mjuk). 
Den hårda latexen användes för att kunna göra tester på prover som ännu inte filmbildat när de torkat vid rumstemperatur och den mjuka latexen användes för att göra referens prover mot bestrykningen med hård latex.
Resultaten visade att det går att mäta styvhetsökning i bestrykningen som en följd av filmformation med DMTA och filmformation av latex i bestrykningen troligtvis beror på både tid, temperatur och provets historia. 
Ett försök att mäta vilken uppehålls tid vid en specifik temperatur som krävs för att filmbildningen skall fulländas genomfördes. 
Dessa försök visade att DMTA:n inte var en lämplig metod för att mäta denna tid då styvheten verkade öka under en längre tid. 
Detta kan bero på att pigment partiklarna packade sig tätare och på så sätt orsakade en ökning av styvheten. 
Därför gjordes ett annat försök som involverar ugns härdning, men på grund av tidsbrist blev det bara en mätserie utförd. 
Den sist nämnda metoden visade dock goda resultat och måste därför bedömas ha en potential.
Metod: 
Empirin samlades in genom en kvalitativ metod bestående av djupintervjuer med konsumenter som köper lågengagemangsprodukten spaghetti.
Teoretiska perspektiv: 
Teorikapitlet strävar efter att ge en bild av några marknadsföringsbegrepp och förpackningen och dess olika element. 
Till sist presenteras två modeller som ligger till grund för undersökningen.
Empirisk analys: 
Empiri består av tolv stycken djupintervjuer med konsumenter som köper spaghetti. 
Dessa har sedan tolkats och analyserats utifrån modellen om köpbeslutsprocessen, som är uppbyggd av teorierna.
Slutsatser: 
Slutsatserna är att faktorn information är av centralbetydelse för konsumenten i sitt köpbeslut och ur den teoretiska grund som finns i uppsatsen, kan inte alla teorier ges riktighet. 
Av undersökningen framkom det också att graden av engagemang i köpbeslutsprocessen har ökat. 
Enligt konsumenterna ska en optimal förpackning vara återförslutningsbar, vara större och ha refill funktion samt ha en tydlig innehållsdeklaration på svenska. 
Resultatet visar att producenterna måste uppdatera sig med dagens trender.
Klimatfrågan har fått stor uppmärksamhet den senaste tiden i och med de klimatförändringar som har börjat ske på jorden. 
Följden av detta är fler naturolyckor där översvämningar är en fara som kommer att öka världen över. 
Idag är inte Sverige ett särskilt översvämningshotat land, men frekvensen bedöms öka även här. 
I Klimat- och sårbarhetsutredningens delbetänkande har undersökningar gjorts över risker och åtgärder för tre sjöar i Sverige, där Vänerområdet anses vara mycket hotat. 
Vänerns normalnivå är idag 44,54 m, men i ett förändrat klimat är den högsta, dimensionerande nivån (10 000-årsnivå) beräknad till 47,4 m. 
Vid denna nivå uppstår konsekvenser för samhället då en stor del bebyggelse, tung industri och jordbruksmark ligger mycket Vänernära. 
Uppsatsen är kvalitativ och baserad på både intervjuer och litteraturstudier. 
I uppsatsen görs en närmare studie av industrier där Akzo Nobel Base Chemicals är ett exempel. 
För övrigt diskuteras olika konsekvenser som finns för samhället och naturen vid en översvämning av industrier (som dock idag är svåra att förutsäga), vilka förslag på förebyggande som finns och om det finns någon lagstiftning som vidrör frågor kring naturrisker gällande industrier.
Karlstad kommun vill att Karlstad ska uppnå 100 000 invånare, mot idag dryga 80 000. 
För att nå dit måste tätortsnära skogar exploateras. 
För att få reda på hur välbesökta de tätortsnära skogarna är i Karlstad, genomfördes i november 2005, februari, maj och augusti-september 2006 en kvantitativ besöksstudie av I2-skogen i nordvästra Karlstad. 
I2-skogen är ett tätortsnära område omgärdat av bostäder åt tre håll. 
I området finns bland annat flera motionsspår, golfbana och skjutbanor. Studien visar att området är välbesökt, ca 180 000 besökare per år. 77 % av besökarna bor i närområdet runt skogen, inom ett avstånd av 500 meter. 
Boendeformerna i området speglar besökarna och deras aktiviteter och I2-skogen kan kallas för en "vardagsskog" med besökare som återkommer flera dagar i veckan. 
Om de tätortsnära skogarna runt Karlstad exploateras enligt kommunens översiktsplan kommer det att påverka invånare som idag bor nära skogsområden till att de får längre avstånd mellan bostaden och skogen. 
Ett längre avstånd kan göra att det tar för lång tid att ta sig till skogsområden, vilket leder till att antal besök minskar. 
När människor inte har tid att vistas i skogen ökar stress och ohälsa, även barn påverkas negativt av att inte få leka fritt i en tätortsnära skog. 
Det är nu läge att inrätta någon form av områdesskydd för vissa av de tätortsnära skogarna runt Karlstad, då de har ett oerhört viktigt socialt värde för befolkningen i Karlstad och därför behöver bevaras för framtiden.
Bakgrund: De svenska börsbolagen gör större vinster än någonsin tidigare, men har fått stor kritik för att vara för långsamma i sin vinstallokering. 
Företag med överkapitaliserade balansräkningar utan investeringsbehov är potentiella måltavlor för riskkapitalisternas affärsidé om finansiell effektivisering och en aggressivare kapitalstruktur. 
Debatten i media har skapat kritik kring dessa så kallade kortsiktiga och giriga bolagsplundrare som påstås förstöra finansiella värden och kreditvärdigheten i företagen. 
I tidigare fall har marknaden svarat positivt på riskkapitalisternas investeringar, något som har reflekterats i ett kraftigt ökande aktiepris. 
Skeptiker hävdar dock att spekulationer är anledningen till att marknadsvärdet drivs upp, inte fundamentala aspekter.
Syfte: 
Syftet med denna magisteruppsats är att fastställa en bild av fenomenet riskkapital och hur dess aktiva ägande inverkar på svenska börsbolags kreditbetyg, kapitalstruktur och värdering.
Metod: 
För att uppnå syftet med vår magisteruppsats har en kvalitativ ansats till-lämpats baserad på tre börsbolag där riskkapitalisters aktiva ägande spelat en betydande roll. 
Det empiriska materialet har insamlats genom personliga intervjuer med aktie- och kreditanalytiker, och studien förlitar sig även på markandsdata, artiklar och nyhetssändningar i media, samt respektive bolags kvartals- och årsrapporter.
Slutsats: Studien har gjorts over den tidsperiod som varit riskkapitalisternas inve-steringshorisont – explicit och implicit. 
Genom att analysera det aktiva ägarskapet i tre svenska börsbolag kan slutsatsen dras att det inverkat positivt i form av högre prestanda och marknadsvärdering. 
De finansiella förändringarna har, till skillnad från kritiken, styrkt kreditbetyget i fallen Lindex och Volvo. 
En analys av Skandia/Old Mutual visade dock en marginellt ökad kreditrisk. 
Slutsatsen visar härmed att riskkapitalisternas inverkan på svenska börsbolag är värdeförädlande utan att äventyra den finansiella statusen.
Sammanfattning
Enligt världshälsoorganisationen WHO:s hälsorapport från 2002 utgör fysisk inaktivitet och fetma tillsammans mer än 10 procent av den globala samlade sjukdomsbördan och ger upphov till ökande kostnader för hälso- och sjukvården. 
WHO bedömer att 80 procent av hjärt-kärlsjukdomarna, 90 procent av diabetes typ 2 och 30 procent av all cancer kan förebyggas genom bra matvanor, tillräckligt med fysisk aktivitet och genom att sluta röka.
Med denna undersökning vill jag undersöka gymnasieelevers kostvanor samt se om det finns skillnader mellan pojkar och flickors kostvanor.
Undersökningen har gjorts med en kvantitativ ansats där gymnasieelever i årskurs ett, två och tre har svarat på frågor i en enkät. 
Svarsalternativen i enkäten var strukturerade så att eleverna fick fylla i ett eller flera alternativ som stämde överens med deras kostvanor. 
Tre frågor hade ett skattningsalternativ.
För att ha en bra kosthållning bör man äta frukost, lunch och middag samt ett till tre mellanmål och att detta fördelas så jämt som möjligt över dagen. 
Man bör också äta rikligt med fullkornprodukter, frukt och grönsaker.
Resultatet visar att de flesta elever äter frukost, lunch och middag men att ett fåtal elever äter mellanmål. 
De flesta elever har en hälsosam kosthållning. 
Flickor äter mer frukt och grönsaker än pojkar. 
Pojkar dricker mer läsk och light läsk samt att pojkar äter mer godis, chips och choklad än flickor.
Slutsatsen är att eleverna överlag äter hälsosamt vilket kan bero på tidningar och TV som ständigt informerar oss om risker med övervikt och fetma. 
Ofta kan vi läsa i tidningar eller se TV om hur vi ska äta för att må bra och gå ner i vikt. 
Det kan vara så att eleverna har kunskap om vad som är hälsosamt men att de ändå inte klarar att motstå frestelsen för godis, chips och choklad. 
Det kan bero på det utbud av godis, chips och choklad som finns lättillgängligt bland annat i affärer, kiosker och bensinmackar. 
En ide om att få eleverna att äta mer frukt är att elevrestaurangen serverar frukt dagligen.
Med anledning av att allt färre elever väljer språk som tillval på gymnasiet så är syftet med detta examensarbete att ta reda på vad som påverkar gymnasieelever att välja, respektive välja bort, språk som tillval. 
Det jag främst vill undersöka är ifall det finns skillnader i motivation, attityder och nöjdhet/missnöje med undervisningen mellan de som har valt språk och de som har valt bort språk som tillval. 
Vidare syftar undersökningen till att ta reda på vilka förbättringar både elever och lärare tycker vore nödvändiga. 
Metoden som användes var både kvalitativ och kvantitativ i form av intervjuer och två olika enkäter. 
Fyra elever och två lärare intervjuades och enkäterna besvarades av 34 elever med språk som tillval och av 40 elever med andra tillval. 
Resultatet visar inte på några specifika skillnader förutom motivation mellan grupperna, däremot fann jag flera möjliga orsaker till bortval; bland annat ointresse, taktikval och tråkig undervisning. 
De förbättringar som efterfrågades var till viss del organisatoriska, men till största delen handlade de om själva undervisningen. 
Det jag kom fram till är att undervisningen på högstadiet troligen påverkar bortvalen i hög grad och att det är förbättringar där, samt ett nytt skolsystem som premierar språk, som är de viktigaste faktorerna för att få fler elever att välja språk som tillval.
Den här rapporten behandlar ett examensarbete i integrerad produktutveckling. Examensarbetet har gjorts i samarbete med företaget Kinnarps AB.
Uppdraget bestod i att utveckla en ny stol till café och lunchrum som ska möta marknadens förväntningar och krav samt passa in i Kinnarps AB:s sortiment. 
Under projektet har det förutom rena konstruktions- och designförslag gjorts alltifrån marknadsanalys för att få reda på marknadens och kundernas krav, kartläggning av och anpassning till produktion och validering med bl a framtagning av prototyp.
Resultatet av arbetet är en stålrörsstol, vars like inte finns i Kinnarps AB:s sortiment idag. 
Stolen har ett underrede i bockat stålrör samt separat sits och rygg, precis som de befintliga stolarna, Jig och Tango, som den är tänkt att ersätta. 
Det som är speciellt med stolen och som urskiljer den från konkurrenternas stolar är den mycket greppvänliga ryggen och den sviktande rörelsen i ryggen. 
Den införda svikten är något nytt för den här typen av stolar och finns idag varken i Kinnarps AB:s sortiment eller ute på marknaden.
Produktutvecklingsprocessen är en iterativ process som kan beskrivas med aktiviteterna: fastställande av kundkrav, kravspecifikation, konceptgenerering, utvärdering, förkroppsligande samt detaljdesign. 
Att veta vad marknaden vill ha eller behöver är en avgörande faktor för en lyckad produkt. 
Marknadsanalysen visade att den nya stolen bör vara en bekväm och inbjudande stol som är lätt och enkel med en tidlös design och organiska former. 
Att stolen ska vara möjlig att stapla, hänga upp och koppla ihop med andra stolar visade sig vara viktigt.
Att stolen har bra ergonomi är viktigt, varför olika forskares verk studerats. 
För att ytterligare undersöka de ergonomiska aspekterna har en analys gjorts i programmet SAMMIE.
För att göra en ordentlig uppföljning och utvärdering av resultatet togs det fram en prototyp. 
Det kommer även att göras en riskanalys och kvalitetstest i Kinnarps AB:s ackrediterade laboratorium.
Förhoppningsvis har arbetet resulterat i en stol med hög kvalitet och som har god potential att synas i konkurrensen på marknaden.
Denna uppsats undersöker vilka faktorer som påverkar förändringar i elspotpriset på Nord Pool. 
Avsikten är att resultatet skall ligga till grund för en prisuppskattningsmodell för Lunds Energikoncernen AB. 
Faktorerna bestämdes genom en förstudie där viktig litteratur om elmarknaden studerades samt samtal med Lunds Energikoncernen AB. 
De faktorer som undersöks i denna uppsats är priset på utsläppsrätter, nettoexport till Tysk-land, temperatur, nederbörd, priset på kol och villaolja samt konjunkturutveckling i Sve-rige.
Undersökningen av faktorerna bestod av en multipel regressionsanalys med undersökta faktorer som oberoende variabler och elspotpriset på Nord Pool som den beroende va-riabeln. 
Faktorerna blev indelade i två grupper dagsgruppen och månadsgruppen, grunden till uppdelningen är som namnen antyder att statistiken var observerad dygnsvis och må-nadsvis. 
I månadsgruppen ingick nettoexport till Tyskland, priset på kol, villaolja samt konjunktur och ur denna grupp visade sig endast nettoexport till Tyskland ha statistisk signifikans.
I dagsgruppen ingick de faktorer som oftast omnämns i litteraturen som prispåverkande, nämligen temperatur, nederbörd och priset på utsläppsrätter. 
Dock visade sig nederbörd inte ha någon statistisk signifikant påverkan på elpriset varvid ett nytt test på ett nytt sta-tistiskt underlag gjordes för nederbörden vilket gav samma resultat, vilket var förvånan-de. 
Både temperatur och priset på utsläppsrätter visade sig dock ha statistisk signifikans och detta intygades genom ytterligare test.
Härefter gjordes en regressionsanalys med de faktorer visat sig ha statistisk signifikans som oberoende variabler, det vill säga nettoexport till Tyskland, temperatur och priset på utsläppsrätter gentemot elpriset som beroende variabel. 
Denna enkla prognosmodell kunde förklara så mycket som 70 procent av förändringarna i elpriset.
Slutligen diskuteras prognosmodellen av författarna, en brist är bland annat att den inte kan förutse hastiga förändringar i priset och att den behöver kalibreras om när den nya handelsperioden för utsläppsrätter sätter i gång 2008. 
Dock gav analysen positiva signa-ler om att det kan vara möjligt att basera en prismodell på el med de faktorer som har störst inverkan på den dyraste produktionsteknologi som oftast används i elproduktio-nen, då elmarknaden i praktiken tillämpar marginalprissättning.
